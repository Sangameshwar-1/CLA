* Test file for 2-input XOR gate (xor22 - Magic extracted)
* ==========================================================

.include "/home/sangam/Documents/VLSI_PROJ_2017/MAGIC/TSMC_180nm.txt"

* SPICE3 file created from xor22.ext - technology: scmos
.option scale=0.09u

.subckt xor2 a0 b0 p0 vdd gnd

* Node mapping from xor22.spice:
* 3 = a0 (input A)
* 6 = b0 (input B)  
* 2 = abar (a0 inverted)
* 5 = bbar (b0 inverted)
* a_59_1237# = b0 connection node
* p0 = output

* SPICE3 file created from xor22.ext - technology: scmos

.option scale=0.09u

M1000 a_164_1182# 3 vdd w_158_1153# CMOSP w=80 l=2
+  ad=480 pd=172 as=880 ps=352
M1001 a_266_1166# 4 p0 Gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=400 ps=180
M1002 p0 3 a_266_1182# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1003 gnd 5 a_266_1166# Gnd CMOSN w=40 l=2
+  ad=440 pd=192 as=0 ps=0
M1004 a_164_1166# 6 p0 w_158_1153# CMOSP w=80 l=2
+  ad=480 pd=172 as=800 ps=340
M1005 vdd 3 5 w_89_1106# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1006 vdd a_59_1237# 4 w_90_1226# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1007 p0 4 a_164_1182# w_158_1153# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 a_266_1182# 6 gnd Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 gnd 3 5 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1010 vdd 4 a_164_1166# w_158_1153# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 gnd a_59_1237# 4 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
C0 gnd a_266_1166# 0.41fF
C1 p0 a_266_1182# 0.45fF
C2 vdd 5 0.84fF
C3 w_158_1153# p0 0.21fF
C4 w_158_1153# 6 0.06fF
C5 4 a_59_1237# 0.05fF
C6 vdd w_89_1106# 0.11fF
C7 p0 a_266_1166# 0.45fF
C8 4 vdd 0.84fF
C9 5 w_89_1106# 0.06fF
C10 4 5 0.07fF
C11 gnd a_59_1237# 0.05fF
C12 w_158_1153# 3 0.08fF
C13 p0 a_164_1166# 0.82fF
C14 gnd vdd 0.40fF
C15 w_158_1153# a_164_1182# 0.01fF
C16 gnd 5 0.21fF
C17 6 a_59_1237# 0.05fF
C18 vdd p0 0.03fF
C19 gnd 4 0.28fF
C20 vdd 6 0.31fF
C21 p0 5 0.04fF
C22 6 5 0.05fF
C23 4 p0 0.17fF
C24 4 6 0.57fF
C25 vdd 3 0.29fF
C26 vdd a_164_1182# 0.86fF
C27 w_90_1226# a_59_1237# 0.06fF
C28 5 3 0.05fF
C29 w_90_1226# vdd 0.11fF
C30 gnd p0 0.03fF
C31 gnd 6 0.73fF
C32 3 w_89_1106# 0.06fF
C33 4 3 1.36fF
C34 w_90_1226# 4 0.06fF
C35 6 p0 0.01fF
C36 gnd 3 0.12fF
C37 w_158_1153# a_164_1166# 0.01fF
C38 p0 3 0.17fF
C39 6 3 0.19fF
C40 w_158_1153# vdd 0.05fF
C41 p0 a_164_1182# 0.82fF
C42 w_158_1153# 4 0.14fF
C43 vdd a_164_1166# 0.82fF
C44 gnd a_266_1182# 0.41fF
C45 vdd a_59_1237# 0.02fF
C46 a_266_1166# Gnd 0.01fF
C47 5 Gnd 1.45fF
C48 a_266_1182# Gnd 0.01fF
C49 6 Gnd 0.06fF
C50 3 Gnd 1.02fF
C51 p0 Gnd 0.28fF
C52 4 Gnd 2.61fF
C53 vdd Gnd 1.72fF
C54 a_59_1237# Gnd 0.15fF
C55 gnd Gnd 5.76fF
C56 w_89_1106# Gnd 1.35fF
C57 w_158_1153# Gnd 4.44fF
C58 w_90_1226# Gnd 1.35fF


.ends xor2

* ========== TESTBENCH ==========

.param SUPPLY=1.8
.global gnd vdd

VDD vdd gnd {SUPPLY}

* Test 1: A0=0, B0=0 -> P0=0
VA_00 a0_00 gnd 0
VB_00 b0_00 gnd 0
Xxor_00 a0_00 b0_00 p0_00 vdd gnd xor2
Cload_00 p0_00 gnd 10f

* Test 2: A0=0, B0=1 -> P0=1
VA_01 a0_01 gnd 0
VB_01 b0_01 gnd {SUPPLY}
Xxor_01 a0_01 b0_01 p0_01 vdd gnd xor2
Cload_01 p0_01 gnd 10f

* Test 3: A0=1, B0=0 -> P0=1
VA_10 a0_10 gnd {SUPPLY}
VB_10 b0_10 gnd 0
Xxor_10 a0_10 b0_10 p0_10 vdd gnd xor2
Cload_10 p0_10 gnd 10f

* Test 4: A0=1, B0=1 -> P0=0
VA_11 a0_11 gnd {SUPPLY}
VB_11 b0_11 gnd {SUPPLY}
Xxor_11 a0_11 b0_11 p0_11 vdd gnd xor2
Cload_11 p0_11 gnd 10f

* Dynamic test
VA_dyn a0_dyn gnd PULSE(0 {SUPPLY} 1n 100p 100p 2n 4n)
VB_dyn b0_dyn gnd PULSE(0 {SUPPLY} 2n 100p 100p 4n 8n)
Xxor_dyn a0_dyn b0_dyn p0_dyn vdd gnd xor2
Cload_dyn p0_dyn gnd 10f

.control
set numdgt=12

echo ""
echo "=========================================="
echo "  2-INPUT XOR GATE TEST (xor22)"
echo "=========================================="
echo "  P0 = A0 XOR B0"
echo ""

op

echo "Truth Table:"
echo "  A0 B0 | P0 | Expected"
echo "  ------+----+---------"

if v(p0_00) < 0.3
  echo "  0  0  | 0  |    0     PASS"
else
  echo "  0  0  | 1  |    0     FAIL"
end

if v(p0_01) > 1.5
  echo "  0  1  | 1  |    1     PASS"
else
  echo "  0  1  | 0  |    1     FAIL"
end

if v(p0_10) > 1.5
  echo "  1  0  | 1  |    1     PASS"
else
  echo "  1  0  | 0  |    1     FAIL"
end

if v(p0_11) < 0.3
  echo "  1  1  | 0  |    0     PASS"
else
  echo "  1  1  | 1  |    0     FAIL"
end

echo ""
echo "Internal Nodes (Test 00: A0=0, B0=0):"
echo "  Node 2 (abar): " v(xxor_00.2) "V"
echo "  Node 5 (bbar): " v(xxor_00.5) "V"
echo "  Node 3 (a0):   " v(xxor_00.3) "V"
echo "  Node 6 (b0):   " v(xxor_00.6) "V"
echo ""

tran 10p 10n

* Plot A0, B0, P0
plot v(a0_dyn) v(b0_dyn)+2 v(p0_dyn)+4 title 'XOR22: Inputs and Output'

* Plot internal nodes 2,3,5,6
plot v(xxor_dyn.2) v(xxor_dyn.3)+2 v(xxor_dyn.5)+4 v(xxor_dyn.6)+6 title 'XOR22: Internal Nodes 2,3,5,6'

* Plot all together
plot v(a0_dyn) v(xxor_dyn.2)+2 v(b0_dyn)+4 v(xxor_dyn.5)+6 v(p0_dyn)+8 title 'XOR22: Complete Signal Set'

.endc
.end