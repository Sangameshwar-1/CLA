magic
tech scmos
timestamp 1763386411
<< nwell >>
rect -11 71 21 163
<< ntransistor >>
rect 0 45 2 55
rect 8 45 10 55
<< ptransistor >>
rect 0 77 2 157
rect 8 77 10 157
<< ndiffusion >>
rect -1 45 0 55
rect 2 45 3 55
rect 7 45 8 55
rect 10 45 11 55
<< pdiffusion >>
rect -1 77 0 157
rect 2 77 3 157
rect 7 77 8 157
rect 10 77 11 157
<< ndcontact >>
rect -5 45 -1 55
rect 3 45 7 55
rect 11 45 15 55
<< pdcontact >>
rect -5 77 -1 157
rect 3 77 7 157
rect 11 77 15 157
<< polysilicon >>
rect 0 157 2 170
rect 8 157 10 170
rect 0 55 2 77
rect 8 55 10 77
rect 0 42 2 45
rect 8 42 10 45
<< polycontact >>
rect -1 170 3 174
rect 7 170 11 174
<< metal1 >>
rect -1 174 3 180
rect 7 174 11 180
rect 11 157 15 166
rect -5 64 -1 77
rect -5 59 15 64
rect -5 55 -1 59
rect 11 55 15 59
rect 3 37 7 45
<< labels >>
rlabel metal1 -5 62 -1 66 1 out
rlabel metal1 -5 63 -1 67 1 nor_2
rlabel metal1 7 176 11 180 5 b
rlabel metal1 -1 176 3 180 5 a
rlabel metal1 11 162 15 166 1 vdd
rlabel metal1 3 37 7 41 1 gnd
<< end >>
