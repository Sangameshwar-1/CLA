* Generate sum outputs (S)
* S_i = P_i XOR C_i
.subckt si p0 p1 p2 p3 p4 c0 c1 c2 c3 c4 s0 s1 s2 s3 s4 vdd gnd 
Xxor0 p0 c0 s0 vdd gnd xor2
Xxor1 p1 c1 s1 vdd gnd xor2
Xxor2 p2 c2 s2 vdd gnd xor2
Xxor3 p3 c3 s3 vdd gnd xor2
Xxor4 p4 c4 s4 vdd gnd xor2
.ends si