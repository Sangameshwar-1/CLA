magic
tech scmos
timestamp 1763529985
<< nwell >>
rect -58 480 -34 536
rect 62 479 86 535
rect -11 375 37 467
<< ntransistor >>
rect -47 544 -45 564
rect 73 543 75 563
rect 0 319 2 359
rect 8 319 10 359
rect 16 319 18 359
rect 24 319 26 359
<< ptransistor >>
rect -47 490 -45 530
rect 73 489 75 529
rect 0 381 2 461
rect 8 381 10 461
rect 16 381 18 461
rect 24 381 26 461
<< ndiffusion >>
rect -48 544 -47 564
rect -45 544 -44 564
rect 72 543 73 563
rect 75 543 76 563
rect -1 319 0 359
rect 2 319 3 359
rect 7 319 8 359
rect 10 319 11 359
rect 15 319 16 359
rect 18 319 19 359
rect 23 319 24 359
rect 26 319 27 359
<< pdiffusion >>
rect -48 490 -47 530
rect -45 490 -44 530
rect 72 489 73 529
rect 75 489 76 529
rect -1 381 0 461
rect 2 381 3 461
rect 7 381 8 461
rect 10 381 11 461
rect 15 381 16 461
rect 18 381 19 461
rect 23 381 24 461
rect 26 381 27 461
<< ndcontact >>
rect -52 544 -48 564
rect -44 544 -40 564
rect 68 543 72 563
rect 76 543 80 563
rect -5 319 -1 359
rect 3 319 7 359
rect 11 319 15 359
rect 19 319 23 359
rect 27 319 31 359
<< pdcontact >>
rect -52 490 -48 530
rect -44 490 -40 530
rect 68 489 72 529
rect 76 489 80 529
rect -5 381 -1 461
rect 3 381 7 461
rect 11 381 15 461
rect 19 381 23 461
rect 27 381 31 461
<< polysilicon >>
rect -47 564 -45 567
rect 73 563 75 566
rect -47 530 -45 544
rect 73 529 75 543
rect -47 487 -45 490
rect 73 486 75 489
rect 0 461 2 474
rect 8 461 10 474
rect 16 461 18 474
rect 24 461 26 474
rect 0 378 2 381
rect 8 370 10 381
rect 0 368 10 370
rect 16 370 18 381
rect 24 378 26 381
rect 16 368 26 370
rect 0 359 2 368
rect 8 359 10 362
rect 16 359 18 362
rect 24 359 26 368
rect 0 316 2 319
rect 8 311 10 319
rect 2 309 10 311
rect 16 311 18 319
rect 24 316 26 319
rect 16 309 25 311
<< polycontact >>
rect -45 537 -41 541
rect 75 536 79 540
rect -1 474 3 478
rect 7 474 11 478
rect 15 474 19 478
rect 23 474 27 478
rect -2 308 2 312
rect 25 308 29 312
<< metal1 >>
rect -75 568 -40 572
rect -75 464 -71 568
rect -44 564 -40 568
rect -52 541 -48 544
rect 15 541 19 597
rect 76 568 80 569
rect 76 564 102 568
rect 76 563 80 564
rect -66 537 -48 541
rect -41 537 19 541
rect 68 540 72 543
rect -65 475 -61 537
rect -52 530 -48 537
rect -15 506 11 510
rect -44 484 -40 490
rect -31 484 -26 485
rect -58 480 -26 484
rect -15 475 -11 506
rect 0 480 3 494
rect -65 471 -11 475
rect -1 478 3 480
rect 7 478 11 506
rect 15 478 19 537
rect 23 536 72 540
rect 79 536 90 540
rect 23 478 27 536
rect 40 530 44 536
rect 68 529 72 536
rect 48 470 52 484
rect 76 483 80 489
rect 98 484 102 564
rect 62 479 89 483
rect 85 470 89 479
rect 112 470 116 578
rect 11 466 116 470
rect -75 460 -28 464
rect 11 461 15 466
rect -5 368 -1 381
rect 27 368 31 381
rect -14 364 31 368
rect -5 359 -1 364
rect 27 359 31 364
rect 11 308 15 319
rect -1 285 2 308
rect 25 304 28 308
rect 40 285 43 403
rect -1 282 43 285
<< m2contact >>
rect -31 485 -25 491
rect -1 494 4 499
rect 39 525 44 530
rect 48 484 54 490
rect 97 478 103 484
rect -28 459 -22 465
rect 40 403 46 409
rect 10 302 16 308
rect 25 299 30 304
<< metal2 >>
rect 90 587 93 595
rect 0 584 93 587
rect 0 499 3 584
rect 40 502 44 525
rect -25 485 48 489
rect 90 459 93 584
rect -28 281 -24 459
rect 60 456 93 459
rect 41 409 44 423
rect 11 281 15 302
rect 26 294 29 299
rect 60 294 63 456
rect 99 448 103 478
rect 26 291 63 294
rect 68 444 103 448
rect -28 280 17 281
rect 68 280 72 444
rect -28 277 72 280
rect 11 276 72 277
rect 67 269 71 276
<< m3contact >>
rect 40 497 45 502
rect 41 423 46 428
<< metal3 >>
rect 41 428 44 497
<< labels >>
rlabel metal2 67 269 71 273 1 gnd
rlabel metal1 15 591 19 596 1 a
rlabel metal1 112 573 116 578 7 vdd
rlabel metal1 -14 364 -10 368 1 xor
rlabel metal2 90 591 93 595 5 b
<< end >>
