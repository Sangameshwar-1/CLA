magic
tech scmos
timestamp 1764432779
<< nwell >>
rect -405 1149 -353 1181
rect -404 1096 -348 1120
rect -395 1014 -343 1046
rect -395 959 -339 983
rect -365 890 -313 922
rect -364 844 -308 868
rect 88 758 140 790
rect 241 692 293 724
rect -870 548 -818 580
rect 89 566 145 590
rect -778 546 -726 548
rect -945 510 -893 542
rect -779 514 -726 546
rect -873 476 -821 508
rect -94 442 -42 521
rect -873 392 -821 424
rect -781 390 -729 392
rect -948 354 -896 386
rect -782 358 -729 390
rect -94 354 -42 412
rect -876 320 -824 352
rect -94 292 -42 342
rect 188 322 240 401
rect 761 299 813 331
rect 853 297 905 299
rect -877 237 -825 269
rect -94 249 -42 281
rect 686 261 738 293
rect 852 265 905 297
rect -785 235 -733 237
rect -952 199 -900 231
rect -786 203 -733 235
rect 758 227 810 259
rect -880 165 -828 197
rect 758 143 810 175
rect 850 141 902 143
rect -880 79 -828 111
rect -788 77 -736 79
rect -94 78 -42 136
rect 683 105 735 137
rect 849 109 902 141
rect -955 41 -903 73
rect -789 45 -736 77
rect -883 7 -831 39
rect -94 16 -42 66
rect 143 15 195 73
rect 755 71 807 103
rect -94 -27 -42 5
rect 754 -12 806 20
rect 846 -14 898 -12
rect 679 -50 731 -18
rect 845 -46 898 -14
rect 751 -84 803 -52
rect -883 -125 -831 -93
rect -791 -127 -739 -125
rect -958 -163 -906 -131
rect -792 -159 -739 -127
rect -886 -197 -834 -165
rect -94 -200 -42 -150
rect 751 -170 803 -138
rect 843 -172 895 -170
rect -94 -250 -42 -218
rect 108 -231 160 -181
rect 676 -208 728 -176
rect 842 -204 895 -172
rect 748 -242 800 -210
rect -93 -393 -41 -361
rect 748 -374 800 -342
rect 840 -376 892 -374
rect 81 -412 133 -380
rect 673 -412 725 -380
rect 839 -408 892 -376
rect 745 -446 797 -414
<< ntransistor >>
rect -337 1168 -297 1170
rect -337 1160 -297 1162
rect -340 1107 -320 1109
rect -327 1033 -287 1035
rect -327 1025 -287 1027
rect -331 970 -311 972
rect -297 909 -257 911
rect -297 901 -257 903
rect -300 855 -280 857
rect 156 777 196 779
rect 156 769 196 771
rect 309 711 349 713
rect 309 703 349 705
rect 153 577 173 579
rect -802 567 -762 569
rect -802 559 -762 561
rect -710 535 -670 537
rect -877 529 -837 531
rect -710 527 -670 529
rect -877 521 -837 523
rect -26 505 74 507
rect -805 495 -765 497
rect -805 487 -765 489
rect -26 487 74 489
rect -26 479 74 481
rect -26 461 74 463
rect -26 453 74 455
rect -805 411 -765 413
rect -805 403 -765 405
rect -26 399 54 401
rect -26 391 54 393
rect 256 385 356 387
rect -713 379 -673 381
rect -880 373 -840 375
rect -713 371 -673 373
rect -26 373 54 375
rect -880 365 -840 367
rect -26 365 54 367
rect 256 367 356 369
rect 256 359 356 361
rect -808 339 -768 341
rect 256 341 356 343
rect -808 331 -768 333
rect 256 333 356 335
rect -26 329 34 331
rect 829 318 869 320
rect -26 311 34 313
rect 829 310 869 312
rect -26 303 34 305
rect 921 286 961 288
rect 754 280 794 282
rect 921 278 961 280
rect 754 272 794 274
rect -26 268 14 270
rect -26 260 14 262
rect -809 256 -769 258
rect -809 248 -769 250
rect 826 246 866 248
rect 826 238 866 240
rect -717 224 -677 226
rect -884 218 -844 220
rect -717 216 -677 218
rect -884 210 -844 212
rect -812 184 -772 186
rect -812 176 -772 178
rect 826 162 866 164
rect 826 154 866 156
rect -26 123 54 125
rect 918 130 958 132
rect 751 124 791 126
rect -26 115 54 117
rect 918 122 958 124
rect 751 116 791 118
rect -812 98 -772 100
rect -26 97 54 99
rect -812 90 -772 92
rect -26 89 54 91
rect 823 90 863 92
rect 823 82 863 84
rect -720 66 -680 68
rect -887 60 -847 62
rect -720 58 -680 60
rect -887 52 -847 54
rect 211 60 291 62
rect -26 53 34 55
rect 211 52 291 54
rect -26 35 34 37
rect -815 26 -775 28
rect 211 34 291 36
rect -26 27 34 29
rect 211 26 291 28
rect -815 18 -775 20
rect 822 7 862 9
rect 822 -1 862 1
rect -26 -8 14 -6
rect -26 -16 14 -14
rect 914 -25 954 -23
rect 747 -31 787 -29
rect 914 -33 954 -31
rect 747 -39 787 -37
rect 819 -65 859 -63
rect 819 -73 859 -71
rect -815 -106 -775 -104
rect -815 -114 -775 -112
rect -723 -138 -683 -136
rect -890 -144 -850 -142
rect -723 -146 -683 -144
rect -890 -152 -850 -150
rect 819 -151 859 -149
rect 819 -159 859 -157
rect -26 -163 34 -161
rect -818 -178 -778 -176
rect -26 -181 34 -179
rect -818 -186 -778 -184
rect -26 -189 34 -187
rect 911 -183 951 -181
rect 744 -189 784 -187
rect 176 -194 236 -192
rect 911 -191 951 -189
rect 744 -197 784 -195
rect 176 -212 236 -210
rect 176 -220 236 -218
rect 816 -223 856 -221
rect -26 -231 14 -229
rect 816 -231 856 -229
rect -26 -239 14 -237
rect 816 -355 856 -353
rect 816 -363 856 -361
rect -25 -374 15 -372
rect -25 -382 15 -380
rect 149 -393 189 -391
rect 908 -387 948 -385
rect 741 -393 781 -391
rect 149 -401 189 -399
rect 908 -395 948 -393
rect 741 -401 781 -399
rect 813 -427 853 -425
rect 813 -435 853 -433
<< ptransistor >>
rect -399 1168 -359 1170
rect -399 1160 -359 1162
rect -394 1107 -354 1109
rect -389 1033 -349 1035
rect -389 1025 -349 1027
rect -385 970 -345 972
rect -359 909 -319 911
rect -359 901 -319 903
rect -354 855 -314 857
rect 94 777 134 779
rect 94 769 134 771
rect 247 711 287 713
rect 247 703 287 705
rect 99 577 139 579
rect -864 567 -824 569
rect -864 559 -824 561
rect -772 535 -732 537
rect -939 529 -899 531
rect -772 527 -732 529
rect -939 521 -899 523
rect -88 505 -48 507
rect -867 495 -827 497
rect -867 487 -827 489
rect -88 487 -48 489
rect -88 479 -48 481
rect -88 461 -48 463
rect -88 453 -48 455
rect -867 411 -827 413
rect -867 403 -827 405
rect -88 399 -48 401
rect -88 391 -48 393
rect 194 385 234 387
rect -775 379 -735 381
rect -942 373 -902 375
rect -775 371 -735 373
rect -88 373 -48 375
rect -942 365 -902 367
rect -88 365 -48 367
rect 194 367 234 369
rect 194 359 234 361
rect -870 339 -830 341
rect 194 341 234 343
rect -870 331 -830 333
rect 194 333 234 335
rect -88 329 -48 331
rect 767 318 807 320
rect -88 311 -48 313
rect 767 310 807 312
rect -88 303 -48 305
rect 859 286 899 288
rect 692 280 732 282
rect 859 278 899 280
rect 692 272 732 274
rect -88 268 -48 270
rect -88 260 -48 262
rect -871 256 -831 258
rect -871 248 -831 250
rect 764 246 804 248
rect 764 238 804 240
rect -779 224 -739 226
rect -946 218 -906 220
rect -779 216 -739 218
rect -946 210 -906 212
rect -874 184 -834 186
rect -874 176 -834 178
rect 764 162 804 164
rect 764 154 804 156
rect -88 123 -48 125
rect 856 130 896 132
rect 689 124 729 126
rect -88 115 -48 117
rect 856 122 896 124
rect 689 116 729 118
rect -874 98 -834 100
rect -88 97 -48 99
rect -874 90 -834 92
rect -88 89 -48 91
rect 761 90 801 92
rect 761 82 801 84
rect -782 66 -742 68
rect -949 60 -909 62
rect -782 58 -742 60
rect -949 52 -909 54
rect 149 60 189 62
rect -88 53 -48 55
rect 149 52 189 54
rect -88 35 -48 37
rect -877 26 -837 28
rect 149 34 189 36
rect -88 27 -48 29
rect 149 26 189 28
rect -877 18 -837 20
rect 760 7 800 9
rect 760 -1 800 1
rect -88 -8 -48 -6
rect -88 -16 -48 -14
rect 852 -25 892 -23
rect 685 -31 725 -29
rect 852 -33 892 -31
rect 685 -39 725 -37
rect 757 -65 797 -63
rect 757 -73 797 -71
rect -877 -106 -837 -104
rect -877 -114 -837 -112
rect -785 -138 -745 -136
rect -952 -144 -912 -142
rect -785 -146 -745 -144
rect -952 -152 -912 -150
rect 757 -151 797 -149
rect 757 -159 797 -157
rect -88 -163 -48 -161
rect -880 -178 -840 -176
rect -88 -181 -48 -179
rect -880 -186 -840 -184
rect -88 -189 -48 -187
rect 849 -183 889 -181
rect 682 -189 722 -187
rect 114 -194 154 -192
rect 849 -191 889 -189
rect 682 -197 722 -195
rect 114 -212 154 -210
rect 114 -220 154 -218
rect 754 -223 794 -221
rect -88 -231 -48 -229
rect 754 -231 794 -229
rect -88 -239 -48 -237
rect 754 -355 794 -353
rect 754 -363 794 -361
rect -87 -374 -47 -372
rect -87 -382 -47 -380
rect 87 -393 127 -391
rect 846 -387 886 -385
rect 679 -393 719 -391
rect 87 -401 127 -399
rect 846 -395 886 -393
rect 679 -401 719 -399
rect 751 -427 791 -425
rect 751 -435 791 -433
<< ndiffusion >>
rect -337 1170 -297 1171
rect -337 1167 -297 1168
rect -337 1162 -297 1163
rect -337 1159 -297 1160
rect -340 1109 -320 1110
rect -340 1106 -320 1107
rect -327 1035 -287 1036
rect -327 1032 -287 1033
rect -327 1027 -287 1028
rect -327 1024 -287 1025
rect -331 972 -311 973
rect -331 969 -311 970
rect -297 911 -257 912
rect -297 908 -257 909
rect -297 903 -257 904
rect -297 900 -257 901
rect -300 857 -280 858
rect -300 854 -280 855
rect 156 779 196 780
rect 156 776 196 777
rect 156 771 196 772
rect 156 768 196 769
rect 309 713 349 714
rect 309 710 349 711
rect 309 705 349 706
rect 309 702 349 703
rect 153 579 173 580
rect 153 576 173 577
rect -802 569 -762 570
rect -802 566 -762 567
rect -802 561 -762 562
rect -802 558 -762 559
rect -710 537 -670 538
rect -877 531 -837 532
rect -877 528 -837 529
rect -710 534 -670 535
rect -710 529 -670 530
rect -877 523 -837 524
rect -710 526 -670 527
rect -877 520 -837 521
rect -26 507 74 508
rect -26 504 74 505
rect -805 497 -765 498
rect -805 494 -765 495
rect -805 489 -765 490
rect -805 486 -765 487
rect -26 489 74 490
rect -26 486 74 487
rect -26 481 74 482
rect -26 478 74 479
rect -26 463 74 464
rect -26 460 74 461
rect -26 455 74 456
rect -26 452 74 453
rect -805 413 -765 414
rect -805 410 -765 411
rect -805 405 -765 406
rect -805 402 -765 403
rect -26 401 54 402
rect -26 398 54 399
rect -26 393 54 394
rect -26 390 54 391
rect 256 387 356 388
rect -713 381 -673 382
rect 256 384 356 385
rect -880 375 -840 376
rect -880 372 -840 373
rect -713 378 -673 379
rect -713 373 -673 374
rect -26 375 54 376
rect -880 367 -840 368
rect -713 370 -673 371
rect -880 364 -840 365
rect -26 372 54 373
rect -26 367 54 368
rect 256 369 356 370
rect -26 364 54 365
rect 256 366 356 367
rect 256 361 356 362
rect 256 358 356 359
rect -808 341 -768 342
rect 256 343 356 344
rect -808 338 -768 339
rect -808 333 -768 334
rect -808 330 -768 331
rect 256 340 356 341
rect 256 335 356 336
rect -26 331 34 332
rect -26 328 34 329
rect 256 332 356 333
rect 829 320 869 321
rect -26 313 34 314
rect -26 310 34 311
rect 829 317 869 318
rect 829 312 869 313
rect -26 305 34 306
rect 829 309 869 310
rect -26 302 34 303
rect 921 288 961 289
rect 754 282 794 283
rect 754 279 794 280
rect 921 285 961 286
rect 921 280 961 281
rect 754 274 794 275
rect 921 277 961 278
rect -26 270 14 271
rect -26 267 14 268
rect 754 271 794 272
rect -26 262 14 263
rect -809 258 -769 259
rect -809 255 -769 256
rect -26 259 14 260
rect -809 250 -769 251
rect -809 247 -769 248
rect 826 248 866 249
rect 826 245 866 246
rect 826 240 866 241
rect 826 237 866 238
rect -717 226 -677 227
rect -884 220 -844 221
rect -884 217 -844 218
rect -717 223 -677 224
rect -717 218 -677 219
rect -884 212 -844 213
rect -717 215 -677 216
rect -884 209 -844 210
rect -812 186 -772 187
rect -812 183 -772 184
rect -812 178 -772 179
rect -812 175 -772 176
rect 826 164 866 165
rect 826 161 866 162
rect 826 156 866 157
rect 826 153 866 154
rect -26 125 54 126
rect 918 132 958 133
rect 751 126 791 127
rect -26 122 54 123
rect -26 117 54 118
rect 751 123 791 124
rect 918 129 958 130
rect 918 124 958 125
rect 751 118 791 119
rect 918 121 958 122
rect -26 114 54 115
rect 751 115 791 116
rect -812 100 -772 101
rect -812 97 -772 98
rect -26 99 54 100
rect -812 92 -772 93
rect -812 89 -772 90
rect -26 96 54 97
rect -26 91 54 92
rect 823 92 863 93
rect -26 88 54 89
rect 823 89 863 90
rect 823 84 863 85
rect 823 81 863 82
rect -720 68 -680 69
rect -887 62 -847 63
rect -887 59 -847 60
rect -720 65 -680 66
rect -720 60 -680 61
rect -887 54 -847 55
rect -720 57 -680 58
rect 211 62 291 63
rect -26 55 34 56
rect -887 51 -847 52
rect -26 52 34 53
rect 211 59 291 60
rect 211 54 291 55
rect 211 51 291 52
rect -26 37 34 38
rect -815 28 -775 29
rect -26 34 34 35
rect 211 36 291 37
rect -26 29 34 30
rect -815 25 -775 26
rect -26 26 34 27
rect 211 33 291 34
rect 211 28 291 29
rect 211 25 291 26
rect -815 20 -775 21
rect -815 17 -775 18
rect 822 9 862 10
rect 822 6 862 7
rect 822 1 862 2
rect -26 -6 14 -5
rect 822 -2 862 -1
rect -26 -9 14 -8
rect -26 -14 14 -13
rect -26 -17 14 -16
rect 914 -23 954 -22
rect 747 -29 787 -28
rect 747 -32 787 -31
rect 914 -26 954 -25
rect 914 -31 954 -30
rect 747 -37 787 -36
rect 914 -34 954 -33
rect 747 -40 787 -39
rect 819 -63 859 -62
rect 819 -66 859 -65
rect 819 -71 859 -70
rect 819 -74 859 -73
rect -815 -104 -775 -103
rect -815 -107 -775 -106
rect -815 -112 -775 -111
rect -815 -115 -775 -114
rect -723 -136 -683 -135
rect -890 -142 -850 -141
rect -890 -145 -850 -144
rect -723 -139 -683 -138
rect -723 -144 -683 -143
rect -890 -150 -850 -149
rect -723 -147 -683 -146
rect 819 -149 859 -148
rect -890 -153 -850 -152
rect 819 -152 859 -151
rect 819 -157 859 -156
rect -26 -161 34 -160
rect -26 -164 34 -163
rect 819 -160 859 -159
rect -818 -176 -778 -175
rect -818 -179 -778 -178
rect -26 -179 34 -178
rect -818 -184 -778 -183
rect -818 -187 -778 -186
rect -26 -182 34 -181
rect -26 -187 34 -186
rect -26 -190 34 -189
rect 911 -181 951 -180
rect 744 -187 784 -186
rect 176 -192 236 -191
rect 176 -195 236 -194
rect 744 -190 784 -189
rect 911 -184 951 -183
rect 911 -189 951 -188
rect 744 -195 784 -194
rect 911 -192 951 -191
rect 744 -198 784 -197
rect 176 -210 236 -209
rect 176 -213 236 -212
rect 176 -218 236 -217
rect 176 -221 236 -220
rect 816 -221 856 -220
rect -26 -229 14 -228
rect -26 -232 14 -231
rect 816 -224 856 -223
rect 816 -229 856 -228
rect 816 -232 856 -231
rect -26 -237 14 -236
rect -26 -240 14 -239
rect 816 -353 856 -352
rect 816 -356 856 -355
rect 816 -361 856 -360
rect 816 -364 856 -363
rect -25 -372 15 -371
rect -25 -375 15 -374
rect -25 -380 15 -379
rect -25 -383 15 -382
rect 149 -391 189 -390
rect 149 -394 189 -393
rect 908 -385 948 -384
rect 741 -391 781 -390
rect 149 -399 189 -398
rect 149 -402 189 -401
rect 741 -394 781 -393
rect 908 -388 948 -387
rect 908 -393 948 -392
rect 741 -399 781 -398
rect 908 -396 948 -395
rect 741 -402 781 -401
rect 813 -425 853 -424
rect 813 -428 853 -427
rect 813 -433 853 -432
rect 813 -436 853 -435
<< pdiffusion >>
rect -399 1170 -359 1171
rect -399 1167 -359 1168
rect -399 1162 -359 1163
rect -399 1159 -359 1160
rect -394 1109 -354 1110
rect -394 1106 -354 1107
rect -389 1035 -349 1036
rect -389 1032 -349 1033
rect -389 1027 -349 1028
rect -389 1024 -349 1025
rect -385 972 -345 973
rect -385 969 -345 970
rect -359 911 -319 912
rect -359 908 -319 909
rect -359 903 -319 904
rect -359 900 -319 901
rect -354 857 -314 858
rect -354 854 -314 855
rect 94 779 134 780
rect 94 776 134 777
rect 94 771 134 772
rect 94 768 134 769
rect 247 713 287 714
rect 247 710 287 711
rect 247 705 287 706
rect 247 702 287 703
rect 99 579 139 580
rect 99 576 139 577
rect -864 569 -824 570
rect -864 566 -824 567
rect -864 561 -824 562
rect -864 558 -824 559
rect -939 531 -899 532
rect -772 537 -732 538
rect -772 534 -732 535
rect -939 528 -899 529
rect -939 523 -899 524
rect -772 529 -732 530
rect -772 526 -732 527
rect -939 520 -899 521
rect -88 507 -48 508
rect -88 504 -48 505
rect -867 497 -827 498
rect -867 494 -827 495
rect -867 489 -827 490
rect -867 486 -827 487
rect -88 489 -48 490
rect -88 486 -48 487
rect -88 481 -48 482
rect -88 478 -48 479
rect -88 463 -48 464
rect -88 460 -48 461
rect -88 455 -48 456
rect -88 452 -48 453
rect -867 413 -827 414
rect -867 410 -827 411
rect -867 405 -827 406
rect -867 402 -827 403
rect -88 401 -48 402
rect -88 398 -48 399
rect -88 393 -48 394
rect -88 390 -48 391
rect -942 375 -902 376
rect -775 381 -735 382
rect 194 387 234 388
rect 194 384 234 385
rect -775 378 -735 379
rect -942 372 -902 373
rect -942 367 -902 368
rect -775 373 -735 374
rect -88 375 -48 376
rect -88 372 -48 373
rect -775 370 -735 371
rect -942 364 -902 365
rect -88 367 -48 368
rect 194 369 234 370
rect 194 366 234 367
rect -88 364 -48 365
rect 194 361 234 362
rect 194 358 234 359
rect -870 341 -830 342
rect 194 343 234 344
rect 194 340 234 341
rect -870 338 -830 339
rect -870 333 -830 334
rect -870 330 -830 331
rect -88 331 -48 332
rect 194 335 234 336
rect 194 332 234 333
rect -88 328 -48 329
rect -88 313 -48 314
rect 767 320 807 321
rect 767 317 807 318
rect -88 310 -48 311
rect -88 305 -48 306
rect 767 312 807 313
rect 767 309 807 310
rect -88 302 -48 303
rect 692 282 732 283
rect 859 288 899 289
rect 859 285 899 286
rect 692 279 732 280
rect -88 270 -48 271
rect 692 274 732 275
rect 859 280 899 281
rect 859 277 899 278
rect 692 271 732 272
rect -88 267 -48 268
rect -871 258 -831 259
rect -88 262 -48 263
rect -88 259 -48 260
rect -871 255 -831 256
rect -871 250 -831 251
rect -871 247 -831 248
rect 764 248 804 249
rect 764 245 804 246
rect 764 240 804 241
rect 764 237 804 238
rect -946 220 -906 221
rect -779 226 -739 227
rect -779 223 -739 224
rect -946 217 -906 218
rect -946 212 -906 213
rect -779 218 -739 219
rect -779 215 -739 216
rect -946 209 -906 210
rect -874 186 -834 187
rect -874 183 -834 184
rect -874 178 -834 179
rect -874 175 -834 176
rect 764 164 804 165
rect 764 161 804 162
rect 764 156 804 157
rect 764 153 804 154
rect -88 125 -48 126
rect 689 126 729 127
rect 856 132 896 133
rect 856 129 896 130
rect 689 123 729 124
rect -88 122 -48 123
rect -88 117 -48 118
rect 689 118 729 119
rect 856 124 896 125
rect 856 121 896 122
rect 689 115 729 116
rect -88 114 -48 115
rect -874 100 -834 101
rect -874 97 -834 98
rect -874 92 -834 93
rect -88 99 -48 100
rect -88 96 -48 97
rect -874 89 -834 90
rect -88 91 -48 92
rect 761 92 801 93
rect 761 89 801 90
rect -88 88 -48 89
rect 761 84 801 85
rect 761 81 801 82
rect -949 62 -909 63
rect -782 68 -742 69
rect -782 65 -742 66
rect -949 59 -909 60
rect -949 54 -909 55
rect -782 60 -742 61
rect -782 57 -742 58
rect -88 55 -48 56
rect 149 62 189 63
rect 149 59 189 60
rect -88 52 -48 53
rect -949 51 -909 52
rect 149 54 189 55
rect 149 51 189 52
rect -88 37 -48 38
rect -88 34 -48 35
rect -877 28 -837 29
rect -88 29 -48 30
rect 149 36 189 37
rect 149 33 189 34
rect -88 26 -48 27
rect -877 25 -837 26
rect -877 20 -837 21
rect 149 28 189 29
rect 149 25 189 26
rect -877 17 -837 18
rect 760 9 800 10
rect 760 6 800 7
rect -88 -6 -48 -5
rect 760 1 800 2
rect 760 -2 800 -1
rect -88 -9 -48 -8
rect -88 -14 -48 -13
rect -88 -17 -48 -16
rect 685 -29 725 -28
rect 852 -23 892 -22
rect 852 -26 892 -25
rect 685 -32 725 -31
rect 685 -37 725 -36
rect 852 -31 892 -30
rect 852 -34 892 -33
rect 685 -40 725 -39
rect 757 -63 797 -62
rect 757 -66 797 -65
rect 757 -71 797 -70
rect 757 -74 797 -73
rect -877 -104 -837 -103
rect -877 -107 -837 -106
rect -877 -112 -837 -111
rect -877 -115 -837 -114
rect -952 -142 -912 -141
rect -785 -136 -745 -135
rect -785 -139 -745 -138
rect -952 -145 -912 -144
rect -952 -150 -912 -149
rect -785 -144 -745 -143
rect -785 -147 -745 -146
rect 757 -149 797 -148
rect 757 -152 797 -151
rect -952 -153 -912 -152
rect -88 -161 -48 -160
rect 757 -157 797 -156
rect 757 -160 797 -159
rect -88 -164 -48 -163
rect -880 -176 -840 -175
rect -880 -179 -840 -178
rect -880 -184 -840 -183
rect -88 -179 -48 -178
rect -88 -182 -48 -181
rect -880 -187 -840 -186
rect -88 -187 -48 -186
rect -88 -190 -48 -189
rect 114 -192 154 -191
rect 682 -187 722 -186
rect 849 -181 889 -180
rect 849 -184 889 -183
rect 682 -190 722 -189
rect 114 -195 154 -194
rect 682 -195 722 -194
rect 849 -189 889 -188
rect 849 -192 889 -191
rect 682 -198 722 -197
rect 114 -210 154 -209
rect 114 -213 154 -212
rect 114 -218 154 -217
rect 114 -221 154 -220
rect -88 -229 -48 -228
rect 754 -221 794 -220
rect 754 -224 794 -223
rect -88 -232 -48 -231
rect -88 -237 -48 -236
rect 754 -229 794 -228
rect 754 -232 794 -231
rect -88 -240 -48 -239
rect 754 -353 794 -352
rect 754 -356 794 -355
rect 754 -361 794 -360
rect 754 -364 794 -363
rect -87 -372 -47 -371
rect -87 -375 -47 -374
rect -87 -380 -47 -379
rect -87 -383 -47 -382
rect 87 -391 127 -390
rect 87 -394 127 -393
rect 87 -399 127 -398
rect 679 -391 719 -390
rect 846 -385 886 -384
rect 846 -388 886 -387
rect 679 -394 719 -393
rect 87 -402 127 -401
rect 679 -399 719 -398
rect 846 -393 886 -392
rect 846 -396 886 -395
rect 679 -402 719 -401
rect 751 -425 791 -424
rect 751 -428 791 -427
rect 751 -433 791 -432
rect 751 -436 791 -435
<< ndcontact >>
rect -337 1171 -297 1175
rect -337 1163 -297 1167
rect -337 1155 -297 1159
rect -340 1110 -320 1114
rect -340 1102 -320 1106
rect -327 1036 -287 1040
rect -327 1028 -287 1032
rect -327 1020 -287 1024
rect -331 973 -311 977
rect -331 965 -311 969
rect -297 912 -257 916
rect -297 904 -257 908
rect -297 896 -257 900
rect -300 858 -280 862
rect -300 850 -280 854
rect 156 780 196 784
rect 156 772 196 776
rect 156 764 196 768
rect 309 714 349 718
rect 309 706 349 710
rect 309 698 349 702
rect 153 580 173 584
rect -802 570 -762 574
rect 153 572 173 576
rect -802 562 -762 566
rect -802 554 -762 558
rect -877 532 -837 536
rect -710 538 -670 542
rect -877 524 -837 528
rect -710 530 -670 534
rect -710 522 -670 526
rect -877 516 -837 520
rect -26 508 74 512
rect -805 498 -765 502
rect -26 500 74 504
rect -805 490 -765 494
rect -26 490 74 494
rect -805 482 -765 486
rect -26 482 74 486
rect -26 474 74 478
rect -26 464 74 468
rect -26 456 74 460
rect -26 448 74 452
rect -805 414 -765 418
rect -805 406 -765 410
rect -805 398 -765 402
rect -26 402 54 406
rect -26 394 54 398
rect -26 386 54 390
rect -880 376 -840 380
rect -713 382 -673 386
rect 256 388 356 392
rect 256 380 356 384
rect -880 368 -840 372
rect -713 374 -673 378
rect -26 376 54 380
rect -713 366 -673 370
rect -26 368 54 372
rect 256 370 356 374
rect -880 360 -840 364
rect -26 360 54 364
rect 256 362 356 366
rect 256 354 356 358
rect -808 342 -768 346
rect 256 344 356 348
rect -808 334 -768 338
rect -808 326 -768 330
rect -26 332 34 336
rect 256 336 356 340
rect 256 328 356 332
rect -26 324 34 328
rect -26 314 34 318
rect 829 321 869 325
rect -26 306 34 310
rect 829 313 869 317
rect 829 305 869 309
rect -26 298 34 302
rect 754 283 794 287
rect 921 289 961 293
rect -26 271 14 275
rect 754 275 794 279
rect 921 281 961 285
rect 921 273 961 277
rect -809 259 -769 263
rect 754 267 794 271
rect -26 263 14 267
rect -26 255 14 259
rect -809 251 -769 255
rect -809 243 -769 247
rect 826 249 866 253
rect 826 241 866 245
rect 826 233 866 237
rect -884 221 -844 225
rect -717 227 -677 231
rect -884 213 -844 217
rect -717 219 -677 223
rect -717 211 -677 215
rect -884 205 -844 209
rect -812 187 -772 191
rect -812 179 -772 183
rect -812 171 -772 175
rect 826 165 866 169
rect 826 157 866 161
rect 826 149 866 153
rect -26 126 54 130
rect 751 127 791 131
rect 918 133 958 137
rect -26 118 54 122
rect 751 119 791 123
rect 918 125 958 129
rect 918 117 958 121
rect -26 110 54 114
rect 751 111 791 115
rect -812 101 -772 105
rect -812 93 -772 97
rect -26 100 54 104
rect -812 85 -772 89
rect -26 92 54 96
rect 823 93 863 97
rect -26 84 54 88
rect 823 85 863 89
rect 823 77 863 81
rect -887 63 -847 67
rect -720 69 -680 73
rect -887 55 -847 59
rect -720 61 -680 65
rect -720 53 -680 57
rect -26 56 34 60
rect 211 63 291 67
rect -887 47 -847 51
rect -26 48 34 52
rect 211 55 291 59
rect 211 47 291 51
rect -26 38 34 42
rect -815 29 -775 33
rect -26 30 34 34
rect 211 37 291 41
rect -815 21 -775 25
rect -26 22 34 26
rect 211 29 291 33
rect 211 21 291 25
rect -815 13 -775 17
rect 822 10 862 14
rect -26 -5 14 -1
rect 822 2 862 6
rect 822 -6 862 -2
rect -26 -13 14 -9
rect -26 -21 14 -17
rect 747 -28 787 -24
rect 914 -22 954 -18
rect 747 -36 787 -32
rect 914 -30 954 -26
rect 914 -38 954 -34
rect 747 -44 787 -40
rect 819 -62 859 -58
rect 819 -70 859 -66
rect 819 -78 859 -74
rect -815 -103 -775 -99
rect -815 -111 -775 -107
rect -815 -119 -775 -115
rect -890 -141 -850 -137
rect -723 -135 -683 -131
rect -890 -149 -850 -145
rect -723 -143 -683 -139
rect -723 -151 -683 -147
rect 819 -148 859 -144
rect -890 -157 -850 -153
rect -26 -160 34 -156
rect 819 -156 859 -152
rect 819 -164 859 -160
rect -26 -168 34 -164
rect -818 -175 -778 -171
rect -818 -183 -778 -179
rect -26 -178 34 -174
rect -818 -191 -778 -187
rect -26 -186 34 -182
rect -26 -194 34 -190
rect 176 -191 236 -187
rect 744 -186 784 -182
rect 911 -180 951 -176
rect 176 -199 236 -195
rect 744 -194 784 -190
rect 911 -188 951 -184
rect 911 -196 951 -192
rect 744 -202 784 -198
rect 176 -209 236 -205
rect 176 -217 236 -213
rect -26 -228 14 -224
rect 176 -225 236 -221
rect 816 -220 856 -216
rect 816 -228 856 -224
rect -26 -236 14 -232
rect 816 -236 856 -232
rect -26 -244 14 -240
rect 816 -352 856 -348
rect 816 -360 856 -356
rect -25 -371 15 -367
rect 816 -368 856 -364
rect -25 -379 15 -375
rect -25 -387 15 -383
rect 149 -390 189 -386
rect 741 -390 781 -386
rect 908 -384 948 -380
rect 149 -398 189 -394
rect 741 -398 781 -394
rect 908 -392 948 -388
rect 908 -400 948 -396
rect 149 -406 189 -402
rect 741 -406 781 -402
rect 813 -424 853 -420
rect 813 -432 853 -428
rect 813 -440 853 -436
<< pdcontact >>
rect -399 1171 -359 1175
rect -399 1163 -359 1167
rect -399 1155 -359 1159
rect -394 1110 -354 1114
rect -394 1102 -354 1106
rect -389 1036 -349 1040
rect -389 1028 -349 1032
rect -389 1020 -349 1024
rect -385 973 -345 977
rect -385 965 -345 969
rect -359 912 -319 916
rect -359 904 -319 908
rect -359 896 -319 900
rect -354 858 -314 862
rect -354 850 -314 854
rect 94 780 134 784
rect 94 772 134 776
rect 94 764 134 768
rect 247 714 287 718
rect 247 706 287 710
rect 247 698 287 702
rect 99 580 139 584
rect -864 570 -824 574
rect 99 572 139 576
rect -864 562 -824 566
rect -864 554 -824 558
rect -772 538 -732 542
rect -939 532 -899 536
rect -772 530 -732 534
rect -939 524 -899 528
rect -772 522 -732 526
rect -939 516 -899 520
rect -88 508 -48 512
rect -867 498 -827 502
rect -88 500 -48 504
rect -867 490 -827 494
rect -88 490 -48 494
rect -867 482 -827 486
rect -88 482 -48 486
rect -88 474 -48 478
rect -88 464 -48 468
rect -88 456 -48 460
rect -88 448 -48 452
rect -867 414 -827 418
rect -867 406 -827 410
rect -867 398 -827 402
rect -88 402 -48 406
rect -88 394 -48 398
rect -88 386 -48 390
rect 194 388 234 392
rect -775 382 -735 386
rect -942 376 -902 380
rect 194 380 234 384
rect -775 374 -735 378
rect -942 368 -902 372
rect -88 376 -48 380
rect -775 366 -735 370
rect -88 368 -48 372
rect -942 360 -902 364
rect 194 370 234 374
rect -88 360 -48 364
rect 194 362 234 366
rect 194 354 234 358
rect -870 342 -830 346
rect 194 344 234 348
rect -870 334 -830 338
rect 194 336 234 340
rect -88 332 -48 336
rect -870 326 -830 330
rect -88 324 -48 328
rect 194 328 234 332
rect 767 321 807 325
rect -88 314 -48 318
rect 767 313 807 317
rect -88 306 -48 310
rect 767 305 807 309
rect -88 298 -48 302
rect 859 289 899 293
rect 692 283 732 287
rect 859 281 899 285
rect 692 275 732 279
rect -88 271 -48 275
rect 859 273 899 277
rect -88 263 -48 267
rect -871 259 -831 263
rect 692 267 732 271
rect -871 251 -831 255
rect -88 255 -48 259
rect 764 249 804 253
rect -871 243 -831 247
rect 764 241 804 245
rect 764 233 804 237
rect -779 227 -739 231
rect -946 221 -906 225
rect -779 219 -739 223
rect -946 213 -906 217
rect -779 211 -739 215
rect -946 205 -906 209
rect -874 187 -834 191
rect -874 179 -834 183
rect -874 171 -834 175
rect 764 165 804 169
rect 764 157 804 161
rect 764 149 804 153
rect 856 133 896 137
rect -88 126 -48 130
rect 689 127 729 131
rect 856 125 896 129
rect -88 118 -48 122
rect 689 119 729 123
rect 856 117 896 121
rect -88 110 -48 114
rect 689 111 729 115
rect -874 101 -834 105
rect -88 100 -48 104
rect -874 93 -834 97
rect -88 92 -48 96
rect -874 85 -834 89
rect 761 93 801 97
rect -88 84 -48 88
rect 761 85 801 89
rect 761 77 801 81
rect -782 69 -742 73
rect -949 63 -909 67
rect -782 61 -742 65
rect -949 55 -909 59
rect 149 63 189 67
rect -782 53 -742 57
rect -88 56 -48 60
rect 149 55 189 59
rect -949 47 -909 51
rect -88 48 -48 52
rect 149 47 189 51
rect -88 38 -48 42
rect 149 37 189 41
rect -877 29 -837 33
rect -88 30 -48 34
rect 149 29 189 33
rect -877 21 -837 25
rect -88 22 -48 26
rect 149 21 189 25
rect -877 13 -837 17
rect 760 10 800 14
rect 760 2 800 6
rect -88 -5 -48 -1
rect 760 -6 800 -2
rect -88 -13 -48 -9
rect -88 -21 -48 -17
rect 852 -22 892 -18
rect 685 -28 725 -24
rect 852 -30 892 -26
rect 685 -36 725 -32
rect 852 -38 892 -34
rect 685 -44 725 -40
rect 757 -62 797 -58
rect 757 -70 797 -66
rect 757 -78 797 -74
rect -877 -103 -837 -99
rect -877 -111 -837 -107
rect -877 -119 -837 -115
rect -785 -135 -745 -131
rect -952 -141 -912 -137
rect -785 -143 -745 -139
rect -952 -149 -912 -145
rect -785 -151 -745 -147
rect 757 -148 797 -144
rect -952 -157 -912 -153
rect 757 -156 797 -152
rect -88 -160 -48 -156
rect -88 -168 -48 -164
rect 757 -164 797 -160
rect -880 -175 -840 -171
rect -88 -178 -48 -174
rect -880 -183 -840 -179
rect 849 -180 889 -176
rect -88 -186 -48 -182
rect -880 -191 -840 -187
rect 682 -186 722 -182
rect -88 -194 -48 -190
rect 114 -191 154 -187
rect 849 -188 889 -184
rect 682 -194 722 -190
rect 114 -199 154 -195
rect 849 -196 889 -192
rect 682 -202 722 -198
rect 114 -209 154 -205
rect 114 -217 154 -213
rect 754 -220 794 -216
rect -88 -228 -48 -224
rect 114 -225 154 -221
rect 754 -228 794 -224
rect -88 -236 -48 -232
rect 754 -236 794 -232
rect -88 -244 -48 -240
rect 754 -352 794 -348
rect 754 -360 794 -356
rect -87 -371 -47 -367
rect 754 -368 794 -364
rect -87 -379 -47 -375
rect -87 -387 -47 -383
rect 846 -384 886 -380
rect 87 -390 127 -386
rect 679 -390 719 -386
rect 87 -398 127 -394
rect 846 -392 886 -388
rect 679 -398 719 -394
rect 87 -406 127 -402
rect 846 -400 886 -396
rect 679 -406 719 -402
rect 751 -424 791 -420
rect 751 -432 791 -428
rect 751 -440 791 -436
<< polysilicon >>
rect -412 1168 -399 1170
rect -359 1168 -337 1170
rect -297 1168 -294 1170
rect -412 1160 -399 1162
rect -359 1160 -337 1162
rect -297 1160 -294 1162
rect -347 1109 -343 1110
rect -397 1107 -394 1109
rect -354 1107 -340 1109
rect -320 1107 -317 1109
rect -402 1033 -389 1035
rect -349 1033 -327 1035
rect -287 1033 -284 1035
rect -402 1025 -389 1027
rect -349 1025 -327 1027
rect -287 1025 -284 1027
rect -338 972 -334 973
rect -388 970 -385 972
rect -345 970 -331 972
rect -311 970 -308 972
rect -372 909 -359 911
rect -319 909 -297 911
rect -257 909 -254 911
rect -372 901 -359 903
rect -319 901 -297 903
rect -257 901 -254 903
rect -307 857 -303 858
rect -357 855 -354 857
rect -314 855 -300 857
rect -280 855 -277 857
rect 81 777 94 779
rect 134 777 156 779
rect 196 777 199 779
rect 81 769 94 771
rect 134 769 156 771
rect 196 769 199 771
rect 234 711 247 713
rect 287 711 309 713
rect 349 711 352 713
rect 234 703 247 705
rect 287 703 309 705
rect 349 703 352 705
rect 146 579 150 580
rect 96 577 99 579
rect 139 577 153 579
rect 173 577 176 579
rect -877 567 -864 569
rect -824 567 -802 569
rect -762 567 -759 569
rect -877 559 -864 561
rect -824 559 -802 561
rect -762 559 -759 561
rect -786 535 -772 537
rect -732 535 -710 537
rect -670 535 -667 537
rect -952 529 -939 531
rect -899 529 -877 531
rect -837 529 -834 531
rect -786 527 -772 529
rect -732 527 -710 529
rect -670 527 -667 529
rect -952 521 -939 523
rect -899 521 -877 523
rect -837 521 -834 523
rect -101 505 -88 507
rect -48 505 -26 507
rect 74 505 77 507
rect -880 495 -867 497
rect -827 495 -805 497
rect -765 495 -762 497
rect -880 487 -867 489
rect -827 487 -805 489
rect -765 487 -762 489
rect -101 487 -88 489
rect -48 487 -26 489
rect 74 487 77 489
rect -101 479 -88 481
rect -48 479 -26 481
rect 74 479 77 481
rect -101 461 -88 463
rect -48 461 -26 463
rect 74 461 77 463
rect -101 453 -88 455
rect -48 453 -26 455
rect 74 453 77 455
rect -880 411 -867 413
rect -827 411 -805 413
rect -765 411 -762 413
rect -880 403 -867 405
rect -827 403 -805 405
rect -765 403 -762 405
rect -101 399 -88 401
rect -48 399 -26 401
rect 54 399 57 401
rect -101 391 -88 393
rect -48 391 -26 393
rect 54 391 57 393
rect 181 385 194 387
rect 234 385 256 387
rect 356 385 359 387
rect -789 379 -775 381
rect -735 379 -713 381
rect -673 379 -670 381
rect -955 373 -942 375
rect -902 373 -880 375
rect -840 373 -837 375
rect -789 371 -775 373
rect -735 371 -713 373
rect -673 371 -670 373
rect -101 373 -88 375
rect -48 373 -26 375
rect 54 373 57 375
rect -955 365 -942 367
rect -902 365 -880 367
rect -840 365 -837 367
rect -101 365 -88 367
rect -48 365 -26 367
rect 54 365 57 367
rect 181 367 194 369
rect 234 367 256 369
rect 356 367 359 369
rect 181 359 194 361
rect 234 359 256 361
rect 356 359 359 361
rect -883 339 -870 341
rect -830 339 -808 341
rect -768 339 -765 341
rect 181 341 194 343
rect 234 341 256 343
rect 356 341 359 343
rect -883 331 -870 333
rect -830 331 -808 333
rect -768 331 -765 333
rect 181 333 194 335
rect 234 333 256 335
rect 356 333 359 335
rect -101 329 -88 331
rect -48 329 -26 331
rect 34 329 37 331
rect 754 318 767 320
rect 807 318 829 320
rect 869 318 872 320
rect -101 311 -88 313
rect -48 311 -26 313
rect 34 311 37 313
rect 754 310 767 312
rect 807 310 829 312
rect 869 310 872 312
rect -101 303 -88 305
rect -48 303 -26 305
rect 34 303 37 305
rect 845 286 859 288
rect 899 286 921 288
rect 961 286 964 288
rect 679 280 692 282
rect 732 280 754 282
rect 794 280 797 282
rect 845 278 859 280
rect 899 278 921 280
rect 961 278 964 280
rect 679 272 692 274
rect 732 272 754 274
rect 794 272 797 274
rect -101 268 -88 270
rect -48 268 -26 270
rect 14 268 17 270
rect -101 260 -88 262
rect -48 260 -26 262
rect 14 260 17 262
rect -884 256 -871 258
rect -831 256 -809 258
rect -769 256 -766 258
rect -884 248 -871 250
rect -831 248 -809 250
rect -769 248 -766 250
rect 751 246 764 248
rect 804 246 826 248
rect 866 246 869 248
rect 751 238 764 240
rect 804 238 826 240
rect 866 238 869 240
rect -793 224 -779 226
rect -739 224 -717 226
rect -677 224 -674 226
rect -959 218 -946 220
rect -906 218 -884 220
rect -844 218 -841 220
rect -793 216 -779 218
rect -739 216 -717 218
rect -677 216 -674 218
rect -959 210 -946 212
rect -906 210 -884 212
rect -844 210 -841 212
rect -887 184 -874 186
rect -834 184 -812 186
rect -772 184 -769 186
rect -887 176 -874 178
rect -834 176 -812 178
rect -772 176 -769 178
rect 751 162 764 164
rect 804 162 826 164
rect 866 162 869 164
rect 751 154 764 156
rect 804 154 826 156
rect 866 154 869 156
rect -101 123 -88 125
rect -48 123 -26 125
rect 54 123 57 125
rect 842 130 856 132
rect 896 130 918 132
rect 958 130 961 132
rect 676 124 689 126
rect 729 124 751 126
rect 791 124 794 126
rect -101 115 -88 117
rect -48 115 -26 117
rect 54 115 57 117
rect 842 122 856 124
rect 896 122 918 124
rect 958 122 961 124
rect 676 116 689 118
rect 729 116 751 118
rect 791 116 794 118
rect -887 98 -874 100
rect -834 98 -812 100
rect -772 98 -769 100
rect -101 97 -88 99
rect -48 97 -26 99
rect 54 97 57 99
rect -887 90 -874 92
rect -834 90 -812 92
rect -772 90 -769 92
rect -101 89 -88 91
rect -48 89 -26 91
rect 54 89 57 91
rect 748 90 761 92
rect 801 90 823 92
rect 863 90 866 92
rect 748 82 761 84
rect 801 82 823 84
rect 863 82 866 84
rect -796 66 -782 68
rect -742 66 -720 68
rect -680 66 -677 68
rect -962 60 -949 62
rect -909 60 -887 62
rect -847 60 -844 62
rect -796 58 -782 60
rect -742 58 -720 60
rect -680 58 -677 60
rect -962 52 -949 54
rect -909 52 -887 54
rect -847 52 -844 54
rect 136 60 149 62
rect 189 60 211 62
rect 291 60 294 62
rect -101 53 -88 55
rect -48 53 -26 55
rect 34 53 37 55
rect 136 52 149 54
rect 189 52 211 54
rect 291 52 294 54
rect -101 35 -88 37
rect -48 35 -26 37
rect 34 35 37 37
rect -890 26 -877 28
rect -837 26 -815 28
rect -775 26 -772 28
rect 136 34 149 36
rect 189 34 211 36
rect 291 34 294 36
rect -101 27 -88 29
rect -48 27 -26 29
rect 34 27 37 29
rect 136 26 149 28
rect 189 26 211 28
rect 291 26 294 28
rect -890 18 -877 20
rect -837 18 -815 20
rect -775 18 -772 20
rect 747 7 760 9
rect 800 7 822 9
rect 862 7 865 9
rect 747 -1 760 1
rect 800 -1 822 1
rect 862 -1 865 1
rect -101 -8 -88 -6
rect -48 -8 -26 -6
rect 14 -8 17 -6
rect -101 -16 -88 -14
rect -48 -16 -26 -14
rect 14 -16 17 -14
rect 838 -25 852 -23
rect 892 -25 914 -23
rect 954 -25 957 -23
rect 672 -31 685 -29
rect 725 -31 747 -29
rect 787 -31 790 -29
rect 838 -33 852 -31
rect 892 -33 914 -31
rect 954 -33 957 -31
rect 672 -39 685 -37
rect 725 -39 747 -37
rect 787 -39 790 -37
rect 744 -65 757 -63
rect 797 -65 819 -63
rect 859 -65 862 -63
rect 744 -73 757 -71
rect 797 -73 819 -71
rect 859 -73 862 -71
rect -890 -106 -877 -104
rect -837 -106 -815 -104
rect -775 -106 -772 -104
rect -890 -114 -877 -112
rect -837 -114 -815 -112
rect -775 -114 -772 -112
rect -799 -138 -785 -136
rect -745 -138 -723 -136
rect -683 -138 -680 -136
rect -965 -144 -952 -142
rect -912 -144 -890 -142
rect -850 -144 -847 -142
rect -799 -146 -785 -144
rect -745 -146 -723 -144
rect -683 -146 -680 -144
rect -965 -152 -952 -150
rect -912 -152 -890 -150
rect -850 -152 -847 -150
rect 744 -151 757 -149
rect 797 -151 819 -149
rect 859 -151 862 -149
rect 744 -159 757 -157
rect 797 -159 819 -157
rect 859 -159 862 -157
rect -101 -163 -88 -161
rect -48 -163 -26 -161
rect 34 -163 37 -161
rect -893 -178 -880 -176
rect -840 -178 -818 -176
rect -778 -178 -775 -176
rect -101 -181 -88 -179
rect -48 -181 -26 -179
rect 34 -181 37 -179
rect -893 -186 -880 -184
rect -840 -186 -818 -184
rect -778 -186 -775 -184
rect -101 -189 -88 -187
rect -48 -189 -26 -187
rect 34 -189 37 -187
rect 835 -183 849 -181
rect 889 -183 911 -181
rect 951 -183 954 -181
rect 669 -189 682 -187
rect 722 -189 744 -187
rect 784 -189 787 -187
rect 101 -194 114 -192
rect 154 -194 176 -192
rect 236 -194 239 -192
rect 835 -191 849 -189
rect 889 -191 911 -189
rect 951 -191 954 -189
rect 669 -197 682 -195
rect 722 -197 744 -195
rect 784 -197 787 -195
rect 101 -212 114 -210
rect 154 -212 176 -210
rect 236 -212 239 -210
rect 101 -220 114 -218
rect 154 -220 176 -218
rect 236 -220 239 -218
rect 741 -223 754 -221
rect 794 -223 816 -221
rect 856 -223 859 -221
rect -101 -231 -88 -229
rect -48 -231 -26 -229
rect 14 -231 17 -229
rect 741 -231 754 -229
rect 794 -231 816 -229
rect 856 -231 859 -229
rect -101 -239 -88 -237
rect -48 -239 -26 -237
rect 14 -239 17 -237
rect 741 -355 754 -353
rect 794 -355 816 -353
rect 856 -355 859 -353
rect 741 -363 754 -361
rect 794 -363 816 -361
rect 856 -363 859 -361
rect -100 -374 -87 -372
rect -47 -374 -25 -372
rect 15 -374 18 -372
rect -100 -382 -87 -380
rect -47 -382 -25 -380
rect 15 -382 18 -380
rect 74 -393 87 -391
rect 127 -393 149 -391
rect 189 -393 192 -391
rect 832 -387 846 -385
rect 886 -387 908 -385
rect 948 -387 951 -385
rect 666 -393 679 -391
rect 719 -393 741 -391
rect 781 -393 784 -391
rect 74 -401 87 -399
rect 127 -401 149 -399
rect 189 -401 192 -399
rect 832 -395 846 -393
rect 886 -395 908 -393
rect 948 -395 951 -393
rect 666 -401 679 -399
rect 719 -401 741 -399
rect 781 -401 784 -399
rect 738 -427 751 -425
rect 791 -427 813 -425
rect 853 -427 856 -425
rect 738 -435 751 -433
rect 791 -435 813 -433
rect 853 -435 856 -433
<< polycontact >>
rect -416 1167 -412 1171
rect -416 1159 -412 1163
rect -347 1110 -343 1114
rect -406 1032 -402 1036
rect -406 1024 -402 1028
rect -338 973 -334 977
rect -376 908 -372 912
rect -376 900 -372 904
rect -307 858 -303 862
rect 77 776 81 780
rect 77 768 81 772
rect 230 710 234 714
rect 230 702 234 706
rect 146 580 150 584
rect -881 566 -877 570
rect -881 558 -877 562
rect -956 528 -952 532
rect -790 534 -786 538
rect -956 520 -952 524
rect -790 526 -786 530
rect -105 504 -101 508
rect -884 494 -880 498
rect -884 486 -880 490
rect -105 486 -101 490
rect -105 478 -101 482
rect -105 460 -101 464
rect -105 452 -101 456
rect -884 410 -880 414
rect -884 402 -880 406
rect -105 398 -101 402
rect -105 390 -101 394
rect -959 372 -955 376
rect -793 378 -789 382
rect 177 384 181 388
rect -959 364 -955 368
rect -793 370 -789 374
rect -105 372 -101 376
rect -105 364 -101 368
rect 177 366 181 370
rect 177 358 181 362
rect -887 338 -883 342
rect 177 340 181 344
rect -887 330 -883 334
rect -105 328 -101 332
rect 177 332 181 336
rect -105 310 -101 314
rect 750 317 754 321
rect -105 302 -101 306
rect 750 309 754 313
rect 675 279 679 283
rect 841 285 845 289
rect -105 267 -101 271
rect 675 271 679 275
rect 841 277 845 281
rect -888 255 -884 259
rect -105 259 -101 263
rect -888 247 -884 251
rect 747 245 751 249
rect 747 237 751 241
rect -963 217 -959 221
rect -797 223 -793 227
rect -963 209 -959 213
rect -797 215 -793 219
rect -891 183 -887 187
rect -891 175 -887 179
rect 747 161 751 165
rect 747 153 751 157
rect -105 122 -101 126
rect 672 123 676 127
rect 838 129 842 133
rect -105 114 -101 118
rect 672 115 676 119
rect 838 121 842 125
rect -891 97 -887 101
rect -891 89 -887 93
rect -105 96 -101 100
rect -105 88 -101 92
rect 744 89 748 93
rect 744 81 748 85
rect -966 59 -962 63
rect -800 65 -796 69
rect -966 51 -962 55
rect -800 57 -796 61
rect -105 52 -101 56
rect 132 59 136 63
rect 132 51 136 55
rect -105 34 -101 38
rect -894 25 -890 29
rect -105 26 -101 30
rect 132 33 136 37
rect -894 17 -890 21
rect 132 25 136 29
rect 743 6 747 10
rect -105 -9 -101 -5
rect 743 -2 747 2
rect -105 -17 -101 -13
rect 668 -32 672 -28
rect 834 -26 838 -22
rect 668 -40 672 -36
rect 834 -34 838 -30
rect 740 -66 744 -62
rect 740 -74 744 -70
rect -894 -107 -890 -103
rect -894 -115 -890 -111
rect -969 -145 -965 -141
rect -803 -139 -799 -135
rect -969 -153 -965 -149
rect -803 -147 -799 -143
rect 740 -152 744 -148
rect -105 -164 -101 -160
rect 740 -160 744 -156
rect -897 -179 -893 -175
rect -897 -187 -893 -183
rect -105 -182 -101 -178
rect -105 -190 -101 -186
rect 97 -195 101 -191
rect 665 -190 669 -186
rect 831 -184 835 -180
rect 665 -198 669 -194
rect 831 -192 835 -188
rect 97 -213 101 -209
rect 97 -221 101 -217
rect -105 -232 -101 -228
rect 737 -224 741 -220
rect -105 -240 -101 -236
rect 737 -232 741 -228
rect 737 -356 741 -352
rect 737 -364 741 -360
rect -104 -375 -100 -371
rect -104 -383 -100 -379
rect 70 -394 74 -390
rect 70 -402 74 -398
rect 662 -394 666 -390
rect 828 -388 832 -384
rect 662 -402 666 -398
rect 828 -396 832 -392
rect 734 -428 738 -424
rect 734 -436 738 -432
<< metal1 >>
rect -408 1193 90 1194
rect -408 1190 762 1193
rect -1100 1167 -416 1171
rect -408 1167 -404 1190
rect 86 1189 762 1190
rect -292 1175 -90 1176
rect -359 1171 -351 1175
rect -297 1172 -90 1175
rect -297 1171 -289 1172
rect -1100 -151 -1096 1167
rect -408 1163 -399 1167
rect -1087 1159 -416 1163
rect -1087 598 -1083 1159
rect -408 1150 -404 1163
rect -355 1159 -351 1171
rect -359 1155 -337 1159
rect -293 1158 -289 1171
rect -347 1153 -342 1155
rect -288 1153 -287 1157
rect -408 1146 -400 1150
rect -404 1114 -400 1146
rect -347 1135 -343 1153
rect -293 1152 -289 1153
rect -348 1131 -343 1135
rect -347 1114 -343 1131
rect -316 1114 -311 1119
rect -404 1110 -394 1114
rect -320 1110 -311 1114
rect -404 1094 -400 1110
rect -354 1102 -340 1106
rect -404 1090 -395 1094
rect -1089 588 -1083 598
rect -1077 1032 -406 1036
rect -399 1032 -395 1090
rect -347 1083 -343 1102
rect -316 1098 -311 1110
rect -316 1094 -280 1098
rect -284 1040 -280 1094
rect -349 1036 -341 1040
rect -287 1036 -273 1040
rect -1089 -140 -1084 588
rect -1077 87 -1073 1032
rect -399 1028 -389 1032
rect -1066 1024 -406 1028
rect -1066 118 -1062 1024
rect -399 1014 -395 1028
rect -345 1024 -341 1036
rect -277 1033 -273 1036
rect -273 1028 -272 1032
rect -349 1020 -327 1024
rect -399 1010 -392 1014
rect -396 983 -392 1010
rect -338 1007 -334 1020
rect -338 1003 -168 1007
rect -396 977 -391 983
rect -338 977 -334 1003
rect -307 977 -303 981
rect -396 973 -385 977
rect -311 973 -303 977
rect -396 959 -391 973
rect -345 965 -331 969
rect -396 956 -392 959
rect -396 952 -365 956
rect -1054 908 -376 912
rect -369 908 -365 952
rect -338 950 -334 965
rect -307 963 -303 973
rect -307 959 -248 963
rect -252 916 -248 959
rect -319 912 -311 916
rect -257 914 -248 916
rect -257 912 -240 914
rect -1054 210 -1050 908
rect -369 904 -359 908
rect -1040 900 -376 904
rect -1040 222 -1036 900
rect -369 889 -365 904
rect -315 900 -311 912
rect -252 910 -240 912
rect -244 906 -240 910
rect -240 901 -239 905
rect -319 896 -297 900
rect -172 897 -168 1003
rect -369 885 -362 889
rect -366 868 -362 885
rect -307 883 -303 896
rect -167 892 -166 896
rect -307 879 -201 883
rect -366 862 -360 868
rect -307 862 -303 879
rect -276 862 -272 864
rect -366 858 -354 862
rect -280 858 -272 862
rect -366 844 -360 858
rect -314 850 -300 854
rect -307 846 -303 850
rect -366 838 -362 844
rect -277 844 -272 858
rect -205 861 -201 879
rect -200 856 -199 860
rect -402 834 -362 838
rect -277 831 -273 844
rect -1028 780 75 784
rect -1028 779 77 780
rect -1028 366 -1023 779
rect 71 776 77 779
rect 86 776 90 1189
rect 200 784 204 1172
rect 134 780 142 784
rect 196 780 204 784
rect 85 772 94 776
rect -1016 768 77 772
rect 85 770 90 772
rect -1016 765 -1012 768
rect -1016 755 -1010 765
rect -1015 377 -1010 755
rect -873 756 -869 757
rect -1002 709 -895 714
rect -1002 522 -997 709
rect -992 700 -901 704
rect -992 533 -988 700
rect -962 566 -881 570
rect -873 566 -869 751
rect -666 574 -662 742
rect 85 599 89 770
rect 138 768 142 780
rect 134 764 156 768
rect 146 608 150 764
rect 200 759 204 780
rect 200 756 399 759
rect 177 755 399 756
rect 177 752 204 755
rect 146 604 162 608
rect 85 595 93 599
rect -824 570 -816 574
rect -762 570 -662 574
rect 89 584 93 595
rect 146 584 150 604
rect 177 584 181 752
rect 214 710 230 714
rect 239 710 243 739
rect 374 736 378 739
rect 395 736 399 755
rect 374 732 399 736
rect 374 718 378 732
rect 287 714 295 718
rect 349 714 378 718
rect 214 709 229 710
rect 238 706 247 710
rect 208 704 230 706
rect 205 702 230 704
rect 205 700 213 702
rect 89 580 99 584
rect 173 580 181 584
rect 89 570 93 580
rect 139 572 153 576
rect -962 534 -958 566
rect -873 562 -864 566
rect -887 558 -881 562
rect -962 533 -957 534
rect -992 532 -957 533
rect -899 532 -891 536
rect -992 529 -956 532
rect -977 528 -956 529
rect -962 527 -957 528
rect -948 524 -939 528
rect -962 522 -956 524
rect -1002 520 -956 522
rect -1002 517 -957 520
rect -961 490 -957 517
rect -948 513 -944 524
rect -895 520 -891 532
rect -886 520 -882 558
rect -873 547 -869 562
rect -820 558 -816 570
rect -824 554 -802 558
rect -813 538 -809 554
rect -666 542 -662 570
rect -837 532 -829 536
rect -813 534 -790 538
rect -782 534 -778 542
rect -732 538 -724 542
rect -670 538 -662 542
rect -833 522 -829 532
rect -782 530 -772 534
rect -813 526 -790 530
rect -899 516 -877 520
rect -890 515 -882 516
rect -890 498 -886 515
rect -890 494 -884 498
rect -876 494 -872 508
rect -827 498 -819 502
rect -876 490 -867 494
rect -961 486 -884 490
rect -965 410 -884 414
rect -876 410 -872 490
rect -823 486 -819 498
rect -813 486 -809 526
rect -782 513 -778 530
rect -728 526 -724 538
rect -732 522 -710 526
rect -720 515 -716 522
rect -765 498 -761 502
rect -666 502 -662 538
rect -97 566 93 570
rect -97 529 -93 566
rect -97 521 -92 529
rect -134 504 -133 508
rect -128 504 -105 508
rect -96 504 -92 521
rect -48 508 -40 512
rect 74 508 99 512
rect -756 498 -662 502
rect -97 500 -88 504
rect -827 482 -805 486
rect -666 460 -662 498
rect -669 455 -662 460
rect -410 464 -406 491
rect -122 486 -105 490
rect -96 486 -92 500
rect -44 494 -40 508
rect -48 490 -40 494
rect -32 500 -26 504
rect -32 494 -28 500
rect 95 498 99 508
rect 146 506 150 572
rect 177 498 181 580
rect 95 494 181 498
rect -32 490 -26 494
rect 95 490 99 494
rect -97 482 -88 486
rect -388 478 -105 482
rect -410 460 -105 464
rect -96 460 -92 482
rect -44 478 -40 490
rect -48 474 -39 478
rect -32 474 -26 478
rect -44 468 -40 474
rect -48 464 -40 468
rect -32 468 -28 474
rect -32 464 -26 468
rect -669 418 -665 455
rect -827 414 -819 418
rect -765 414 -665 418
rect -965 378 -961 410
rect -876 406 -867 410
rect -890 402 -884 406
rect -965 377 -960 378
rect -1015 376 -960 377
rect -902 376 -894 380
rect -1015 372 -959 376
rect -965 371 -960 372
rect -951 368 -942 372
rect -965 366 -959 368
rect -1028 364 -959 366
rect -1028 361 -960 364
rect -964 334 -960 361
rect -951 357 -947 368
rect -898 364 -894 376
rect -889 364 -885 402
rect -876 391 -872 406
rect -823 402 -819 414
rect -827 398 -805 402
rect -816 382 -812 398
rect -669 386 -665 414
rect -840 376 -832 380
rect -816 378 -793 382
rect -785 378 -781 386
rect -735 382 -727 386
rect -673 382 -665 386
rect -836 366 -832 376
rect -785 374 -775 378
rect -816 370 -793 374
rect -902 360 -880 364
rect -893 359 -885 360
rect -893 342 -889 359
rect -893 338 -887 342
rect -879 338 -875 352
rect -830 342 -822 346
rect -879 334 -870 338
rect -964 330 -887 334
rect -879 284 -875 334
rect -826 330 -822 342
rect -816 330 -812 370
rect -785 357 -781 374
rect -731 370 -727 382
rect -735 366 -713 370
rect -723 359 -719 366
rect -768 342 -764 346
rect -669 346 -665 382
rect -759 342 -665 346
rect -830 326 -808 330
rect -669 305 -665 342
rect -880 279 -875 284
rect -673 299 -665 305
rect -673 291 -669 299
rect -673 279 -668 291
rect -969 255 -888 259
rect -880 255 -876 279
rect -673 263 -669 279
rect -831 259 -823 263
rect -769 259 -669 263
rect -969 223 -965 255
rect -880 251 -871 255
rect -894 247 -888 251
rect -969 222 -964 223
rect -1040 221 -964 222
rect -906 221 -898 225
rect -1040 218 -963 221
rect -982 217 -963 218
rect -969 216 -964 217
rect -955 213 -946 217
rect -969 211 -963 213
rect -980 210 -963 211
rect -1054 209 -963 210
rect -1054 206 -964 209
rect -968 179 -964 206
rect -955 202 -951 213
rect -902 209 -898 221
rect -893 209 -889 247
rect -880 236 -876 251
rect -827 247 -823 259
rect -831 243 -809 247
rect -820 227 -816 243
rect -673 231 -669 259
rect -844 221 -836 225
rect -820 223 -797 227
rect -789 223 -785 231
rect -739 227 -731 231
rect -677 227 -669 231
rect -840 211 -836 221
rect -789 219 -779 223
rect -820 215 -797 219
rect -906 205 -884 209
rect -897 204 -889 205
rect -897 187 -893 204
rect -897 183 -891 187
rect -883 183 -879 197
rect -834 187 -826 191
rect -883 179 -874 183
rect -968 175 -891 179
rect -1077 82 -1071 87
rect -1066 86 -1059 118
rect -1076 53 -1071 82
rect -1064 64 -1059 86
rect -972 97 -891 101
rect -883 97 -879 179
rect -830 175 -826 187
rect -820 175 -816 215
rect -789 202 -785 219
rect -735 215 -731 227
rect -739 211 -717 215
rect -727 204 -723 211
rect -772 187 -768 191
rect -673 191 -669 227
rect -763 187 -669 191
rect -834 171 -812 175
rect -673 150 -669 187
rect -676 144 -669 150
rect -676 105 -672 144
rect -834 101 -826 105
rect -772 101 -672 105
rect -972 65 -968 97
rect -883 93 -874 97
rect -897 89 -891 93
rect -972 64 -967 65
rect -1064 63 -967 64
rect -909 63 -901 67
rect -1064 59 -966 63
rect -972 58 -967 59
rect -958 55 -949 59
rect -972 53 -966 55
rect -1076 51 -966 53
rect -1076 48 -967 51
rect -971 21 -967 48
rect -958 44 -954 55
rect -905 51 -901 63
rect -896 51 -892 89
rect -883 78 -879 93
rect -830 89 -826 101
rect -834 85 -812 89
rect -823 69 -819 85
rect -676 73 -672 101
rect -847 63 -839 67
rect -823 65 -800 69
rect -792 65 -788 73
rect -742 69 -734 73
rect -680 69 -672 73
rect -843 53 -839 63
rect -792 61 -782 65
rect -823 57 -800 61
rect -909 47 -887 51
rect -900 46 -892 47
rect -900 29 -896 46
rect -900 25 -894 29
rect -886 25 -882 39
rect -837 29 -829 33
rect -886 21 -877 25
rect -971 17 -894 21
rect -975 -107 -894 -103
rect -886 -107 -882 21
rect -833 17 -829 29
rect -823 17 -819 57
rect -792 44 -788 61
rect -738 57 -734 69
rect -742 53 -720 57
rect -730 46 -726 53
rect -775 29 -771 33
rect -676 33 -672 69
rect -766 29 -672 33
rect -837 13 -815 17
rect -676 -68 -672 29
rect -410 100 -406 460
rect -97 456 -88 460
rect -118 452 -105 456
rect -135 398 -105 402
rect -96 398 -92 456
rect -44 452 -40 464
rect -48 448 -26 452
rect -36 436 -32 448
rect -36 432 171 436
rect -48 402 -40 406
rect 54 402 95 406
rect -97 394 -88 398
rect -125 390 -105 394
rect -384 372 -105 376
rect -96 372 -92 394
rect -44 390 -40 402
rect -48 386 -39 390
rect -32 386 -26 390
rect 167 388 171 432
rect 239 428 243 706
rect 291 702 295 714
rect 287 698 309 702
rect 298 485 302 698
rect 374 685 378 714
rect 184 424 243 428
rect 184 401 187 424
rect -44 380 -40 386
rect -48 376 -40 380
rect -32 380 -28 386
rect 167 384 177 388
rect 184 384 188 401
rect 395 392 399 732
rect 234 388 242 392
rect 356 388 399 392
rect 416 632 662 636
rect 167 383 171 384
rect 184 380 194 384
rect -32 376 -26 380
rect -97 368 -88 372
rect -118 364 -105 368
rect -96 336 -92 368
rect -44 364 -40 376
rect 79 366 177 370
rect 184 366 188 380
rect 238 374 242 388
rect 234 370 242 374
rect 250 380 256 384
rect 250 374 254 380
rect 250 370 256 374
rect -48 360 -26 364
rect -36 355 -32 360
rect 79 355 83 366
rect 184 362 194 366
rect -36 351 83 355
rect 98 358 177 362
rect -97 332 -88 336
rect 34 332 74 336
rect -130 328 -105 332
rect -127 310 -105 314
rect -96 310 -92 332
rect -48 324 -40 328
rect -44 318 -40 324
rect -48 314 -40 318
rect -32 324 -26 328
rect -32 318 -28 324
rect -32 314 -26 318
rect -97 306 -88 310
rect -118 302 -105 306
rect -122 267 -105 271
rect -96 267 -92 306
rect -44 302 -40 314
rect -48 298 -26 302
rect -33 293 -29 298
rect 98 293 102 358
rect -33 289 102 293
rect 111 340 177 344
rect 184 340 188 362
rect 238 358 242 370
rect 234 354 243 358
rect 250 354 256 358
rect 238 348 242 354
rect 234 344 242 348
rect 250 348 254 354
rect 250 344 256 348
rect -48 271 -40 275
rect 14 271 74 275
rect -97 263 -88 267
rect -151 259 -105 263
rect -151 217 -147 259
rect -96 235 -92 263
rect -44 259 -40 271
rect -48 255 -26 259
rect -33 250 -29 255
rect 111 250 115 340
rect 184 336 194 340
rect 167 332 177 336
rect -33 246 115 250
rect 184 235 188 336
rect 238 332 242 344
rect 394 334 398 388
rect 234 328 256 332
rect 246 286 250 328
rect 416 286 420 632
rect 669 317 750 321
rect 758 317 762 1189
rect 965 325 969 1173
rect 807 321 815 325
rect 869 321 969 325
rect 246 282 421 286
rect 669 285 673 317
rect 758 313 767 317
rect 744 309 750 313
rect 669 284 674 285
rect 448 283 674 284
rect 732 283 740 287
rect -96 231 188 235
rect 448 279 675 283
rect -141 122 -105 126
rect -96 122 -92 231
rect 74 130 78 223
rect 448 138 453 279
rect 669 278 674 279
rect 683 275 692 279
rect 669 273 675 275
rect 494 271 675 273
rect 494 268 674 271
rect 670 241 674 268
rect 683 264 687 275
rect 736 271 740 283
rect 745 271 749 309
rect 758 298 762 313
rect 811 309 815 321
rect 807 305 829 309
rect 818 289 822 305
rect 965 293 969 321
rect 794 283 802 287
rect 818 285 841 289
rect 849 285 853 293
rect 899 289 907 293
rect 961 289 969 293
rect 798 273 802 283
rect 849 281 859 285
rect 818 277 841 281
rect 732 267 754 271
rect 741 266 749 267
rect 741 249 745 266
rect 741 245 747 249
rect 755 245 759 259
rect 804 249 812 253
rect 755 241 764 245
rect 670 237 747 241
rect -48 126 -40 130
rect 54 126 78 130
rect -97 118 -88 122
rect -388 114 -105 118
rect -410 96 -105 100
rect -96 96 -92 118
rect -44 114 -40 126
rect -48 110 -39 114
rect -32 110 -26 114
rect -44 104 -40 110
rect -48 100 -40 104
rect -32 104 -28 110
rect -32 100 -26 104
rect -680 -72 -672 -68
rect -679 -73 -672 -72
rect -497 23 -492 24
rect -679 -99 -675 -73
rect -837 -103 -829 -99
rect -775 -103 -675 -99
rect -975 -139 -971 -107
rect -886 -111 -877 -107
rect -900 -115 -894 -111
rect -987 -140 -982 -139
rect -975 -140 -970 -139
rect -1089 -141 -970 -140
rect -912 -141 -904 -137
rect -1089 -145 -969 -141
rect -975 -146 -970 -145
rect -961 -149 -952 -145
rect -975 -151 -969 -149
rect -1100 -153 -969 -151
rect -1099 -156 -970 -153
rect -974 -183 -970 -156
rect -961 -160 -957 -149
rect -908 -153 -904 -141
rect -899 -153 -895 -115
rect -886 -126 -882 -111
rect -833 -115 -829 -103
rect -837 -119 -815 -115
rect -826 -135 -822 -119
rect -679 -131 -675 -103
rect -850 -141 -842 -137
rect -826 -139 -803 -135
rect -795 -139 -791 -131
rect -745 -135 -737 -131
rect -683 -135 -675 -131
rect -846 -151 -842 -141
rect -795 -143 -785 -139
rect -826 -147 -803 -143
rect -912 -157 -890 -153
rect -903 -158 -895 -157
rect -903 -175 -899 -158
rect -903 -179 -897 -175
rect -889 -179 -885 -165
rect -840 -175 -832 -171
rect -889 -183 -880 -179
rect -974 -187 -897 -183
rect -889 -247 -885 -183
rect -836 -187 -832 -175
rect -826 -187 -822 -147
rect -795 -160 -791 -143
rect -741 -147 -737 -135
rect -745 -151 -723 -147
rect -733 -158 -729 -151
rect -778 -175 -774 -171
rect -679 -171 -675 -135
rect -769 -175 -675 -171
rect -840 -191 -818 -187
rect -679 -215 -675 -175
rect -679 -247 -673 -215
rect -678 -570 -673 -247
rect -497 -481 -492 18
rect -410 23 -406 96
rect -97 92 -88 96
rect -121 88 -105 92
rect -96 60 -92 92
rect -44 88 -40 100
rect -48 84 -26 88
rect 74 85 78 126
rect 407 133 453 138
rect 666 161 747 165
rect 755 161 759 241
rect 808 237 812 249
rect 818 237 822 277
rect 849 264 853 281
rect 903 277 907 289
rect 899 273 921 277
rect 911 266 915 273
rect 866 249 870 253
rect 965 253 969 289
rect 875 249 969 253
rect 804 233 826 237
rect 965 211 969 249
rect 962 206 969 211
rect 962 169 966 206
rect 804 165 812 169
rect 866 165 966 169
rect -36 71 -32 84
rect -36 67 66 71
rect 62 63 66 67
rect -97 56 -88 60
rect 34 56 49 60
rect 62 59 132 63
rect 140 59 144 73
rect 189 63 197 67
rect 291 63 395 67
rect -135 52 -105 56
rect -388 34 -105 38
rect -96 34 -92 56
rect 140 55 149 59
rect -48 48 -40 52
rect -44 42 -40 48
rect -48 38 -40 42
rect -32 48 -26 52
rect 59 51 132 55
rect -32 42 -28 48
rect -32 38 -26 42
rect -97 30 -88 34
rect -120 26 -105 30
rect -410 -178 -406 18
rect -133 -9 -105 -5
rect -96 -9 -92 30
rect -44 26 -40 38
rect -48 22 -26 26
rect -34 18 -30 22
rect 59 18 63 51
rect -34 14 63 18
rect 73 33 132 37
rect 140 33 144 55
rect 193 51 197 63
rect 189 47 198 51
rect 205 47 211 51
rect 193 41 197 47
rect 189 37 197 41
rect 205 41 209 47
rect 205 37 211 41
rect -48 -5 -40 -1
rect 14 -5 49 -1
rect -97 -13 -88 -9
rect -146 -17 -105 -13
rect -96 -46 -92 -13
rect -44 -17 -40 -5
rect -48 -21 -26 -17
rect -37 -25 -33 -21
rect 73 -25 77 33
rect 140 29 149 33
rect 94 25 132 29
rect -37 -29 77 -25
rect 140 -46 144 29
rect 193 25 197 37
rect 189 21 211 25
rect 198 -27 202 21
rect 407 -27 412 133
rect 666 129 670 161
rect 755 157 764 161
rect 741 153 747 157
rect 666 128 671 129
rect 436 126 516 128
rect 537 127 671 128
rect 729 127 737 131
rect 537 126 672 127
rect 436 123 672 126
rect 436 -10 441 123
rect 521 122 526 123
rect 666 122 671 123
rect 680 119 689 123
rect 666 117 672 119
rect 526 115 672 117
rect 526 112 671 115
rect 667 85 671 112
rect 680 108 684 119
rect 733 115 737 127
rect 742 115 746 153
rect 755 142 759 157
rect 808 153 812 165
rect 804 149 826 153
rect 815 133 819 149
rect 962 137 966 165
rect 791 127 799 131
rect 815 129 838 133
rect 846 129 850 137
rect 896 133 904 137
rect 958 133 966 137
rect 795 117 799 127
rect 846 125 856 129
rect 815 121 838 125
rect 729 111 751 115
rect 738 110 746 111
rect 738 93 742 110
rect 738 89 744 93
rect 752 89 756 103
rect 801 93 809 97
rect 752 85 761 89
rect 667 81 744 85
rect 752 35 756 85
rect 805 81 809 93
rect 815 81 819 121
rect 846 108 850 125
rect 900 121 904 133
rect 896 117 918 121
rect 908 110 912 117
rect 863 93 867 97
rect 962 97 966 133
rect 872 93 966 97
rect 801 77 823 81
rect 962 56 966 93
rect 751 30 756 35
rect 958 50 966 56
rect 958 42 962 50
rect 958 30 963 42
rect 198 -31 412 -27
rect 396 -32 412 -31
rect 424 -15 441 -10
rect 662 6 743 10
rect 751 6 755 30
rect 958 14 962 30
rect 800 10 808 14
rect 862 10 962 14
rect -96 -50 144 -46
rect -96 -156 -92 -50
rect 49 -113 53 -69
rect 53 -118 54 -113
rect 49 -120 53 -118
rect -97 -160 -88 -156
rect 34 -160 49 -156
rect -388 -164 -105 -160
rect -410 -182 -105 -178
rect -96 -182 -92 -160
rect -48 -168 -40 -164
rect -44 -174 -40 -168
rect -48 -178 -40 -174
rect -32 -168 -26 -164
rect -32 -174 -28 -168
rect -32 -178 -26 -174
rect -410 -371 -406 -182
rect -124 -190 -122 -186
rect -97 -186 -88 -182
rect -117 -190 -105 -186
rect -394 -232 -393 -228
rect -388 -232 -105 -228
rect -96 -232 -92 -186
rect -44 -190 -40 -178
rect 104 -187 108 -175
rect -48 -194 -26 -190
rect 104 -191 114 -187
rect 236 -191 394 -187
rect -36 -202 -32 -194
rect 60 -195 97 -191
rect 60 -202 64 -195
rect -36 -206 64 -202
rect 72 -213 97 -209
rect 104 -213 108 -191
rect 154 -199 162 -195
rect 158 -205 162 -199
rect 154 -209 162 -205
rect 170 -199 176 -195
rect 170 -205 174 -199
rect 170 -209 176 -205
rect -48 -228 -40 -224
rect 14 -228 49 -224
rect -97 -236 -88 -232
rect -135 -240 -105 -236
rect -96 -265 -92 -236
rect -44 -240 -40 -228
rect -48 -244 -26 -240
rect -35 -249 -31 -244
rect 72 -249 76 -213
rect 104 -217 114 -213
rect 86 -221 97 -217
rect -35 -253 76 -249
rect 104 -265 108 -217
rect 158 -221 162 -209
rect 154 -225 176 -221
rect 166 -247 170 -225
rect 166 -248 278 -247
rect 424 -248 429 -15
rect 662 -26 666 6
rect 751 2 760 6
rect 737 -2 743 2
rect 662 -27 667 -26
rect 166 -251 429 -248
rect 267 -253 429 -251
rect 438 -28 667 -27
rect 725 -28 733 -24
rect 438 -32 668 -28
rect -96 -269 108 -265
rect -410 -375 -104 -371
rect -96 -375 -92 -269
rect 49 -367 53 -279
rect 104 -350 108 -269
rect -47 -371 -39 -367
rect 15 -371 53 -367
rect 79 -354 108 -350
rect -96 -379 -87 -375
rect -118 -383 -104 -379
rect -116 -457 -112 -383
rect -96 -393 -92 -379
rect -43 -383 -39 -371
rect -47 -387 -25 -383
rect -34 -390 -30 -387
rect -34 -394 70 -390
rect 79 -394 83 -354
rect 127 -390 135 -386
rect 189 -390 393 -386
rect 78 -398 87 -394
rect 69 -402 70 -398
rect 79 -400 83 -398
rect 131 -402 135 -390
rect 127 -406 149 -402
rect 138 -419 142 -406
rect 138 -420 256 -419
rect 438 -420 443 -32
rect 662 -33 667 -32
rect 676 -36 685 -32
rect 662 -38 668 -36
rect 470 -40 668 -38
rect 470 -43 667 -40
rect 470 -48 475 -43
rect 663 -70 667 -43
rect 676 -47 680 -36
rect 729 -40 733 -28
rect 738 -40 742 -2
rect 751 -13 755 2
rect 804 -2 808 10
rect 800 -6 822 -2
rect 811 -22 815 -6
rect 958 -18 962 10
rect 787 -28 795 -24
rect 811 -26 834 -22
rect 842 -26 846 -18
rect 892 -22 900 -18
rect 954 -22 962 -18
rect 791 -38 795 -28
rect 842 -30 852 -26
rect 811 -34 834 -30
rect 725 -44 747 -40
rect 734 -45 742 -44
rect 734 -62 738 -45
rect 734 -66 740 -62
rect 748 -66 752 -52
rect 797 -62 805 -58
rect 748 -70 757 -66
rect 663 -74 740 -70
rect 659 -152 740 -148
rect 748 -152 752 -70
rect 801 -74 805 -62
rect 811 -74 815 -34
rect 842 -47 846 -30
rect 896 -34 900 -22
rect 892 -38 914 -34
rect 904 -45 908 -38
rect 859 -62 863 -58
rect 958 -58 962 -22
rect 868 -62 962 -58
rect 797 -78 819 -74
rect 958 -99 962 -62
rect 955 -105 962 -99
rect 955 -144 959 -105
rect 797 -148 805 -144
rect 859 -148 959 -144
rect 659 -184 663 -152
rect 748 -156 757 -152
rect 734 -160 740 -156
rect 659 -185 664 -184
rect 452 -186 664 -185
rect 722 -186 730 -182
rect 452 -190 665 -186
rect 452 -420 457 -190
rect 659 -191 664 -190
rect 673 -194 682 -190
rect 659 -196 665 -194
rect 138 -423 443 -420
rect 246 -425 443 -423
rect 450 -425 457 -420
rect 484 -198 665 -196
rect 484 -201 664 -198
rect 438 -428 443 -425
rect 452 -457 456 -425
rect -116 -461 456 -457
rect 484 -481 489 -201
rect 660 -228 664 -201
rect 673 -205 677 -194
rect 726 -198 730 -186
rect 735 -198 739 -160
rect 748 -171 752 -156
rect 801 -160 805 -148
rect 797 -164 819 -160
rect 808 -180 812 -164
rect 955 -176 959 -148
rect 784 -186 792 -182
rect 808 -184 831 -180
rect 839 -184 843 -176
rect 889 -180 897 -176
rect 951 -180 959 -176
rect 788 -196 792 -186
rect 839 -188 849 -184
rect 808 -192 831 -188
rect 722 -202 744 -198
rect 731 -203 739 -202
rect 731 -220 735 -203
rect 731 -224 737 -220
rect 745 -224 749 -210
rect 794 -220 802 -216
rect 745 -228 754 -224
rect 660 -232 737 -228
rect 656 -356 737 -352
rect 745 -356 749 -228
rect 798 -232 802 -220
rect 808 -232 812 -192
rect 839 -205 843 -188
rect 893 -192 897 -180
rect 889 -196 911 -192
rect 901 -203 905 -196
rect 856 -220 860 -216
rect 955 -216 959 -180
rect 865 -220 959 -216
rect 794 -236 816 -232
rect 955 -317 959 -220
rect 951 -321 959 -317
rect 952 -322 959 -321
rect 952 -348 956 -322
rect 794 -352 802 -348
rect 856 -352 956 -348
rect 656 -388 660 -356
rect 745 -360 754 -356
rect 731 -364 737 -360
rect 656 -389 661 -388
rect -497 -486 489 -481
rect 593 -390 661 -389
rect 719 -390 727 -386
rect 593 -394 662 -390
rect 593 -570 598 -394
rect 656 -395 661 -394
rect 670 -398 679 -394
rect 656 -400 662 -398
rect 612 -402 662 -400
rect 612 -405 661 -402
rect 612 -407 617 -405
rect 657 -432 661 -405
rect 670 -409 674 -398
rect 723 -402 727 -390
rect 732 -402 736 -364
rect 745 -375 749 -360
rect 798 -364 802 -352
rect 794 -368 816 -364
rect 805 -384 809 -368
rect 952 -380 956 -352
rect 781 -390 789 -386
rect 805 -388 828 -384
rect 836 -388 840 -380
rect 886 -384 894 -380
rect 948 -384 956 -380
rect 785 -400 789 -390
rect 836 -392 846 -388
rect 805 -396 828 -392
rect 719 -406 741 -402
rect 728 -407 736 -406
rect 728 -424 732 -407
rect 728 -428 734 -424
rect 742 -428 746 -414
rect 791 -424 799 -420
rect 742 -432 751 -428
rect 657 -436 734 -432
rect 742 -484 746 -432
rect 795 -436 799 -424
rect 805 -436 809 -396
rect 836 -409 840 -392
rect 890 -396 894 -384
rect 886 -400 908 -396
rect 898 -407 902 -400
rect 853 -424 857 -420
rect 952 -420 956 -384
rect 862 -424 956 -420
rect 791 -440 813 -436
rect 952 -467 956 -424
rect -678 -575 598 -570
<< m2contact >>
rect -90 1172 -85 1177
rect -293 1153 -288 1158
rect -316 1119 -311 1124
rect -347 1077 -342 1083
rect -278 1028 -273 1033
rect -307 981 -302 986
rect -338 944 -333 950
rect -245 901 -240 906
rect -172 892 -167 897
rect -276 864 -271 869
rect -407 834 -402 839
rect -307 840 -302 846
rect -205 856 -200 861
rect -277 826 -272 831
rect 199 1172 204 1177
rect -873 751 -868 756
rect -895 709 -890 714
rect -901 700 -896 705
rect -666 742 -661 747
rect 162 604 167 609
rect 209 709 214 714
rect 200 700 205 705
rect -873 542 -868 547
rect -783 542 -778 547
rect -833 517 -828 522
rect -948 508 -943 513
rect -876 508 -871 513
rect -783 508 -778 513
rect -720 510 -715 515
rect -761 498 -756 503
rect -133 504 -128 509
rect -127 486 -122 491
rect 146 501 151 506
rect -393 478 -388 483
rect 95 485 100 490
rect -876 386 -871 391
rect -786 386 -781 391
rect -836 361 -831 366
rect -951 352 -946 357
rect -879 352 -874 357
rect -786 352 -781 357
rect -723 354 -718 359
rect -764 342 -759 347
rect -880 231 -875 236
rect -790 231 -785 236
rect -840 206 -835 211
rect -955 197 -950 202
rect -883 197 -878 202
rect -790 197 -785 202
rect -727 199 -722 204
rect -768 187 -763 192
rect -883 73 -878 78
rect -793 73 -788 78
rect -843 48 -838 53
rect -958 39 -953 44
rect -886 39 -881 44
rect -793 39 -788 44
rect -730 41 -725 46
rect -771 29 -766 34
rect -123 452 -118 457
rect -140 398 -135 403
rect 95 402 100 407
rect -130 390 -125 395
rect -389 372 -384 377
rect 298 480 303 485
rect 662 632 667 637
rect -123 363 -118 368
rect -135 328 -130 333
rect 74 332 79 337
rect -132 310 -127 315
rect -123 302 -118 307
rect -127 267 -122 272
rect 74 271 79 276
rect -152 212 -147 217
rect 162 331 167 336
rect 394 329 399 334
rect 965 1173 970 1178
rect -146 122 -141 127
rect 74 223 79 228
rect 489 268 494 273
rect 758 293 763 298
rect 848 293 853 298
rect 798 268 803 273
rect 683 259 688 264
rect 755 259 760 264
rect -393 114 -388 119
rect -497 18 -492 23
rect -886 -131 -881 -126
rect -796 -131 -791 -126
rect -846 -156 -841 -151
rect -961 -165 -956 -160
rect -889 -165 -884 -160
rect -796 -165 -791 -160
rect -733 -163 -728 -158
rect -774 -175 -769 -170
rect -126 88 -121 93
rect 848 259 853 264
rect 911 261 916 266
rect 870 249 875 254
rect 74 80 79 85
rect -140 52 -135 57
rect 49 56 54 61
rect -393 33 -388 38
rect -125 26 -120 31
rect -410 18 -405 23
rect -138 -9 -133 -4
rect 395 62 400 67
rect 49 -5 54 0
rect -151 -18 -146 -13
rect 89 24 94 29
rect 521 112 526 117
rect 755 137 760 142
rect 845 137 850 142
rect 795 112 800 117
rect 680 103 685 108
rect 752 103 757 108
rect 845 103 850 108
rect 908 105 913 110
rect 867 93 872 98
rect 49 -69 54 -64
rect 48 -118 53 -113
rect -393 -164 -388 -159
rect 49 -160 55 -155
rect -122 -190 -117 -185
rect -393 -232 -388 -227
rect 394 -191 399 -186
rect 49 -228 54 -223
rect -140 -240 -135 -235
rect 81 -222 86 -217
rect 49 -279 54 -274
rect -123 -383 -118 -378
rect 393 -390 398 -385
rect 64 -402 69 -397
rect 470 -53 475 -48
rect 751 -18 756 -13
rect 841 -18 846 -13
rect 791 -43 796 -38
rect 676 -52 681 -47
rect 748 -52 753 -47
rect 841 -52 846 -47
rect 904 -50 909 -45
rect 863 -62 868 -57
rect 748 -176 753 -171
rect 838 -176 843 -171
rect 788 -201 793 -196
rect 673 -210 678 -205
rect 745 -210 750 -205
rect 838 -210 843 -205
rect 901 -208 906 -203
rect 860 -220 865 -215
rect 612 -412 617 -407
rect 745 -380 750 -375
rect 835 -380 840 -375
rect 785 -405 790 -400
rect 670 -414 675 -409
rect 742 -414 747 -409
rect 835 -414 840 -409
rect 898 -412 903 -407
rect 857 -424 862 -419
<< metal2 >>
rect 180 1176 199 1177
rect -85 1172 199 1176
rect 204 1173 965 1177
rect -317 1119 -316 1123
rect -293 1123 -289 1153
rect -311 1119 -289 1123
rect -317 1115 -313 1119
rect -348 1077 -347 1081
rect -346 1037 -342 1077
rect -308 981 -307 985
rect -277 985 -273 1028
rect -227 1016 -222 1021
rect -302 981 -273 985
rect -338 922 -334 944
rect -338 914 -334 917
rect -277 864 -276 868
rect -244 868 -240 901
rect -271 864 -240 868
rect -873 834 -407 838
rect -873 756 -869 834
rect -307 833 -303 840
rect -205 827 -201 856
rect -172 850 -168 892
rect -277 762 -273 826
rect -666 758 -273 762
rect -666 747 -662 758
rect -890 709 209 714
rect -896 700 200 704
rect 167 604 209 608
rect -868 542 -783 547
rect -828 517 -758 520
rect -943 508 -876 513
rect -871 508 -783 513
rect -761 503 -758 517
rect -720 491 -716 510
rect -353 504 -133 508
rect -720 487 -550 491
rect -371 486 -127 490
rect -871 386 -786 391
rect -831 361 -761 364
rect -946 352 -879 357
rect -874 352 -786 357
rect -764 347 -761 361
rect -723 335 -719 354
rect -648 335 -618 336
rect -723 331 -624 335
rect -619 331 -618 335
rect -875 231 -790 236
rect -835 206 -765 209
rect -950 197 -883 202
rect -878 197 -790 202
rect -768 192 -765 206
rect -727 180 -723 199
rect -652 180 -647 181
rect -393 180 -389 478
rect -341 452 -123 456
rect 95 407 99 485
rect 146 473 150 501
rect 125 469 150 473
rect -353 398 -140 402
rect -371 390 -130 394
rect 95 383 99 402
rect 74 379 99 383
rect -332 364 -123 368
rect 74 337 78 379
rect -353 328 -135 332
rect -371 310 -132 314
rect -302 302 -123 306
rect 74 276 78 332
rect -353 267 -127 271
rect 74 228 78 271
rect 125 217 129 469
rect 205 458 209 604
rect -147 213 129 217
rect 135 454 209 458
rect 135 209 139 454
rect 298 444 302 480
rect 146 440 302 444
rect 146 336 150 440
rect 146 332 162 336
rect 161 331 162 332
rect 91 205 139 209
rect 91 190 95 205
rect -727 176 -389 180
rect -878 73 -793 78
rect -485 70 -481 176
rect -393 119 -389 176
rect 90 166 95 190
rect -371 122 -146 126
rect -838 48 -768 51
rect -953 39 -886 44
rect -881 39 -793 44
rect -771 34 -768 48
rect -730 22 -726 41
rect -393 38 -389 114
rect -341 88 -126 92
rect 49 80 74 84
rect 49 61 53 80
rect -371 52 -140 56
rect -655 22 -650 23
rect -730 18 -497 22
rect -492 18 -410 22
rect -881 -131 -796 -126
rect -841 -156 -771 -153
rect -956 -165 -889 -160
rect -884 -165 -796 -160
rect -774 -170 -771 -156
rect -393 -159 -389 33
rect -332 26 -125 30
rect 49 0 53 56
rect 90 29 94 166
rect 88 24 89 28
rect 394 67 398 329
rect 488 273 493 1074
rect 488 268 489 273
rect 488 265 493 268
rect 521 117 526 1071
rect 667 632 1092 636
rect 763 293 848 298
rect 803 268 873 271
rect 688 259 755 264
rect 760 259 848 264
rect 870 254 873 268
rect 911 242 915 261
rect 986 242 991 243
rect 911 238 991 242
rect 760 137 845 142
rect 800 112 870 115
rect 521 111 526 112
rect 685 103 752 108
rect 757 103 845 108
rect 867 98 870 112
rect 908 86 912 105
rect 983 86 988 87
rect 908 82 988 86
rect 394 62 395 67
rect -371 -9 -138 -5
rect -302 -17 -151 -13
rect -162 -23 -158 -17
rect 49 -64 53 -5
rect -200 -91 85 -87
rect 49 -155 53 -118
rect -733 -182 -729 -163
rect 48 -160 49 -158
rect 48 -161 54 -160
rect -658 -182 -615 -181
rect -733 -186 -615 -182
rect -620 -580 -615 -186
rect -393 -227 -389 -164
rect -341 -190 -122 -186
rect 49 -223 53 -161
rect 81 -217 85 -91
rect 394 -186 398 62
rect 756 -18 841 -13
rect 796 -43 866 -40
rect 470 -48 474 -47
rect 681 -52 748 -47
rect 753 -52 841 -47
rect 80 -222 81 -218
rect -393 -233 -389 -232
rect -332 -240 -140 -236
rect -150 -246 -146 -240
rect 49 -274 53 -228
rect -173 -297 -171 -294
rect -166 -297 68 -294
rect -173 -298 68 -297
rect -342 -383 -123 -379
rect 64 -397 68 -298
rect 394 -385 398 -191
rect 394 -392 398 -390
rect 470 -469 474 -53
rect 863 -57 866 -43
rect 904 -69 908 -50
rect 979 -69 984 -68
rect 904 -73 984 -69
rect 753 -176 838 -171
rect 793 -201 863 -198
rect 678 -210 745 -205
rect 750 -210 838 -205
rect 860 -215 863 -201
rect 901 -227 905 -208
rect 976 -227 981 -226
rect 901 -231 981 -227
rect 750 -380 835 -375
rect 613 -407 618 -404
rect 790 -405 860 -402
rect 617 -412 618 -407
rect -479 -473 474 -469
rect 613 -580 618 -412
rect 675 -414 742 -409
rect 747 -414 835 -409
rect 857 -419 860 -405
rect 898 -431 902 -412
rect 973 -431 978 -430
rect 898 -435 978 -431
rect -620 -585 618 -580
<< m3contact >>
rect 488 1074 493 1079
rect -346 1032 -341 1037
rect -338 917 -333 922
rect -307 828 -302 833
rect -172 845 -167 850
rect -205 822 -200 827
rect -358 504 -353 509
rect -550 487 -545 492
rect -376 486 -371 491
rect -624 330 -619 335
rect -346 452 -341 457
rect -358 398 -353 403
rect -376 390 -371 395
rect -337 363 -332 368
rect -358 328 -353 333
rect -376 310 -371 315
rect -307 301 -302 306
rect -358 267 -353 272
rect -376 122 -371 127
rect -485 64 -480 70
rect -346 88 -341 93
rect -376 52 -371 57
rect -337 26 -332 31
rect 521 1071 526 1076
rect -376 -9 -371 -4
rect -307 -18 -302 -13
rect -205 -91 -200 -86
rect -346 -190 -341 -185
rect -337 -240 -332 -235
rect -171 -297 -166 -292
rect -347 -383 -342 -378
rect -484 -473 -479 -468
<< metal3 >>
rect -565 1238 526 1243
rect -565 517 -560 1238
rect -568 512 -560 517
rect -624 336 -617 337
rect -565 336 -560 512
rect -544 1211 493 1216
rect -544 493 -539 1211
rect 488 1080 493 1211
rect 487 1079 494 1080
rect 487 1074 488 1079
rect 493 1074 494 1079
rect 521 1077 526 1238
rect 487 1073 494 1074
rect 520 1076 527 1077
rect 520 1071 521 1076
rect 526 1071 527 1076
rect 520 1070 527 1071
rect -551 492 -539 493
rect -439 525 -353 530
rect -439 492 -434 525
rect -358 509 -353 525
rect -551 487 -550 492
rect -545 487 -434 492
rect -376 491 -371 496
rect -551 486 -544 487
rect -376 395 -371 486
rect -376 336 -371 390
rect -629 335 -371 336
rect -629 331 -624 335
rect -619 331 -371 335
rect -619 330 -617 331
rect -376 315 -371 331
rect -376 127 -371 310
rect -358 403 -353 504
rect -358 333 -353 398
rect -358 272 -353 328
rect -346 457 -343 1032
rect -486 70 -479 71
rect -486 64 -485 70
rect -480 64 -479 70
rect -484 -468 -480 64
rect -376 57 -371 122
rect -376 -4 -371 52
rect -376 -10 -371 -9
rect -346 93 -343 452
rect -337 368 -334 917
rect -173 850 -166 851
rect -173 845 -172 850
rect -167 845 -166 850
rect -173 844 -166 845
rect -307 827 -302 828
rect -206 827 -199 828
rect -346 -185 -343 88
rect -337 31 -334 363
rect -307 306 -304 827
rect -206 822 -205 827
rect -200 822 -199 827
rect -206 821 -199 822
rect -346 -378 -343 -190
rect -337 -235 -334 26
rect -307 -13 -304 301
rect -307 -24 -304 -18
rect -204 -86 -200 821
rect -204 -92 -201 -91
rect -337 -245 -334 -240
rect -171 -292 -167 844
rect -171 -298 -167 -297
rect -346 -384 -343 -383
<< labels >>
rlabel metal1 -992 -145 -987 -140 3 a0
rlabel metal1 -990 -156 -985 -151 3 b0
rlabel metal1 -989 59 -984 64 1 a1
rlabel metal1 -889 -235 -885 -231 1 vdd
rlabel metal1 -679 -218 -675 -214 1 gnd
rlabel metal1 -987 48 -982 53 1 b1
rlabel space -984 206 -979 211 1 b2
rlabel metal1 -980 361 -975 366 1 b3
rlabel metal1 -982 372 -977 377 1 a3
rlabel metal1 -977 517 -972 522 1 b4
rlabel space -979 528 -974 533 1 a4
rlabel space -986 218 -981 223 1 a2
rlabel metal2 1088 632 1092 636 7 cout
rlabel metal2 983 82 987 86 1 s3
rlabel metal2 986 238 990 242 1 s4
rlabel metal2 979 -73 983 -69 1 s2
rlabel metal2 976 -231 980 -227 1 s1
rlabel metal2 973 -435 977 -431 1 s0
rlabel metal2 -720 487 -716 491 1 p4
rlabel space -723 330 -719 334 1 p3
rlabel metal2 -727 176 -723 180 1 p2
rlabel metal2 -730 18 -726 22 1 p1
rlabel metal2 -733 -186 -729 -182 1 p0
rlabel metal2 -338 929 -334 933 1 g1
rlabel metal2 -346 1058 -342 1062 1 g0
rlabel metal3 -307 808 -304 812 1 g2
rlabel metal1 146 527 149 531 1 g3
rlabel space 297 574 300 578 1 g4bar
rlabel metal1 357 -31 360 -27 1 c4
rlabel metal1 347 -253 350 -249 1 c3
rlabel metal1 347 -425 350 -421 1 c2
rlabel metal1 349 -461 352 -457 1 c1
rlabel metal1 380 -575 383 -571 1 c0
<< end >>
