magic
tech scmos
timestamp 1763483110
<< nwell >>
rect -11 71 47 123
<< ntransistor >>
rect 0 -25 2 55
rect 8 -25 10 55
rect 26 -25 28 55
rect 34 -25 36 55
<< ptransistor >>
rect 0 77 2 117
rect 8 77 10 117
rect 26 77 28 117
rect 34 77 36 117
<< ndiffusion >>
rect -1 -25 0 55
rect 2 -25 3 55
rect 7 -25 8 55
rect 10 -25 11 55
rect 25 -25 26 55
rect 28 -25 29 55
rect 33 -25 34 55
rect 36 -25 37 55
<< pdiffusion >>
rect -1 77 0 117
rect 2 77 3 117
rect 7 77 8 117
rect 10 77 11 117
rect 25 77 26 117
rect 28 77 29 117
rect 33 77 34 117
rect 36 77 37 117
<< ndcontact >>
rect -5 -25 -1 55
rect 3 -25 7 55
rect 11 -25 15 55
rect 21 -25 25 55
rect 29 -25 33 55
rect 37 -25 41 55
<< pdcontact >>
rect -5 77 -1 117
rect 3 77 7 117
rect 11 77 15 117
rect 21 77 25 117
rect 29 77 33 117
rect 37 77 41 117
<< polysilicon >>
rect 0 117 2 130
rect 8 117 10 130
rect 26 117 28 130
rect 34 117 36 130
rect 0 55 2 77
rect 8 55 10 77
rect 26 55 28 77
rect 34 55 36 77
rect 0 -28 2 -25
rect 8 -28 10 -25
rect 26 -28 28 -25
rect 34 -28 36 -25
<< polycontact >>
rect -1 130 3 134
rect 7 130 11 134
rect 25 130 29 134
rect 33 130 37 134
<< metal1 >>
rect -1 134 3 140
rect 7 134 11 140
rect 25 134 29 140
rect 33 134 37 140
rect 3 123 33 126
rect 3 117 7 123
rect 29 117 33 123
rect -5 73 -1 77
rect 11 73 15 77
rect 21 73 25 77
rect 37 73 41 77
rect -5 69 41 73
rect -5 55 -1 69
rect 21 68 25 69
rect 11 57 25 61
rect 11 55 15 57
rect 21 55 25 57
rect 37 -33 41 -25
<< labels >>
rlabel metal1 7 136 11 140 5 b
rlabel metal1 -1 136 3 140 5 a
rlabel metal1 -5 62 -1 66 1 out
rlabel metal1 29 122 33 126 1 vdd
rlabel metal1 37 -33 41 -29 1 gnd
rlabel metal1 25 136 29 140 5 c
rlabel metal1 33 136 37 140 5 d
<< end >>
