magic
tech scmos
timestamp 1763562428
<< nwell >>
rect 39 865 91 944
rect 39 777 91 835
rect 39 715 91 765
rect 321 745 373 824
rect 39 672 91 704
rect 39 501 91 559
rect 39 439 91 489
rect 276 438 328 496
rect 39 396 91 428
rect 39 223 91 273
rect 39 173 91 205
rect 241 192 293 242
rect 40 30 92 62
rect 214 11 266 43
<< ntransistor >>
rect 107 928 207 930
rect 107 910 207 912
rect 107 902 207 904
rect 107 884 207 886
rect 107 876 207 878
rect 107 822 187 824
rect 107 814 187 816
rect 389 808 489 810
rect 107 796 187 798
rect 107 788 187 790
rect 389 790 489 792
rect 389 782 489 784
rect 389 764 489 766
rect 389 756 489 758
rect 107 752 167 754
rect 107 734 167 736
rect 107 726 167 728
rect 107 691 147 693
rect 107 683 147 685
rect 107 546 187 548
rect 107 538 187 540
rect 107 520 187 522
rect 107 512 187 514
rect 344 483 424 485
rect 107 476 167 478
rect 344 475 424 477
rect 107 458 167 460
rect 344 457 424 459
rect 107 450 167 452
rect 344 449 424 451
rect 107 415 147 417
rect 107 407 147 409
rect 107 260 167 262
rect 107 242 167 244
rect 107 234 167 236
rect 309 229 369 231
rect 309 211 369 213
rect 309 203 369 205
rect 107 192 147 194
rect 107 184 147 186
rect 108 49 148 51
rect 108 41 148 43
rect 282 30 322 32
rect 282 22 322 24
<< ptransistor >>
rect 45 928 85 930
rect 45 910 85 912
rect 45 902 85 904
rect 45 884 85 886
rect 45 876 85 878
rect 45 822 85 824
rect 45 814 85 816
rect 327 808 367 810
rect 45 796 85 798
rect 45 788 85 790
rect 327 790 367 792
rect 327 782 367 784
rect 327 764 367 766
rect 327 756 367 758
rect 45 752 85 754
rect 45 734 85 736
rect 45 726 85 728
rect 45 691 85 693
rect 45 683 85 685
rect 45 546 85 548
rect 45 538 85 540
rect 45 520 85 522
rect 45 512 85 514
rect 282 483 322 485
rect 45 476 85 478
rect 282 475 322 477
rect 45 458 85 460
rect 282 457 322 459
rect 45 450 85 452
rect 282 449 322 451
rect 45 415 85 417
rect 45 407 85 409
rect 45 260 85 262
rect 45 242 85 244
rect 45 234 85 236
rect 247 229 287 231
rect 247 211 287 213
rect 247 203 287 205
rect 45 192 85 194
rect 45 184 85 186
rect 46 49 86 51
rect 46 41 86 43
rect 220 30 260 32
rect 220 22 260 24
<< ndiffusion >>
rect 107 930 207 931
rect 107 927 207 928
rect 107 912 207 913
rect 107 909 207 910
rect 107 904 207 905
rect 107 901 207 902
rect 107 886 207 887
rect 107 883 207 884
rect 107 878 207 879
rect 107 875 207 876
rect 107 824 187 825
rect 107 821 187 822
rect 107 816 187 817
rect 107 813 187 814
rect 389 810 489 811
rect 389 807 489 808
rect 107 798 187 799
rect 107 795 187 796
rect 107 790 187 791
rect 389 792 489 793
rect 107 787 187 788
rect 389 789 489 790
rect 389 784 489 785
rect 389 781 489 782
rect 389 766 489 767
rect 389 763 489 764
rect 389 758 489 759
rect 107 754 167 755
rect 107 751 167 752
rect 389 755 489 756
rect 107 736 167 737
rect 107 733 167 734
rect 107 728 167 729
rect 107 725 167 726
rect 107 693 147 694
rect 107 690 147 691
rect 107 685 147 686
rect 107 682 147 683
rect 107 548 187 549
rect 107 545 187 546
rect 107 540 187 541
rect 107 537 187 538
rect 107 522 187 523
rect 107 519 187 520
rect 107 514 187 515
rect 107 511 187 512
rect 344 485 424 486
rect 107 478 167 479
rect 107 475 167 476
rect 344 482 424 483
rect 344 477 424 478
rect 344 474 424 475
rect 107 460 167 461
rect 107 457 167 458
rect 344 459 424 460
rect 107 452 167 453
rect 107 449 167 450
rect 344 456 424 457
rect 344 451 424 452
rect 344 448 424 449
rect 107 417 147 418
rect 107 414 147 415
rect 107 409 147 410
rect 107 406 147 407
rect 107 262 167 263
rect 107 259 167 260
rect 107 244 167 245
rect 107 241 167 242
rect 107 236 167 237
rect 107 233 167 234
rect 309 231 369 232
rect 309 228 369 229
rect 309 213 369 214
rect 309 210 369 211
rect 309 205 369 206
rect 309 202 369 203
rect 107 194 147 195
rect 107 191 147 192
rect 107 186 147 187
rect 107 183 147 184
rect 108 51 148 52
rect 108 48 148 49
rect 108 43 148 44
rect 108 40 148 41
rect 282 32 322 33
rect 282 29 322 30
rect 282 24 322 25
rect 282 21 322 22
<< pdiffusion >>
rect 45 930 85 931
rect 45 927 85 928
rect 45 912 85 913
rect 45 909 85 910
rect 45 904 85 905
rect 45 901 85 902
rect 45 886 85 887
rect 45 883 85 884
rect 45 878 85 879
rect 45 875 85 876
rect 45 824 85 825
rect 45 821 85 822
rect 45 816 85 817
rect 45 813 85 814
rect 327 810 367 811
rect 327 807 367 808
rect 45 798 85 799
rect 45 795 85 796
rect 45 790 85 791
rect 327 792 367 793
rect 327 789 367 790
rect 45 787 85 788
rect 327 784 367 785
rect 327 781 367 782
rect 327 766 367 767
rect 327 763 367 764
rect 45 754 85 755
rect 327 758 367 759
rect 327 755 367 756
rect 45 751 85 752
rect 45 736 85 737
rect 45 733 85 734
rect 45 728 85 729
rect 45 725 85 726
rect 45 693 85 694
rect 45 690 85 691
rect 45 685 85 686
rect 45 682 85 683
rect 45 548 85 549
rect 45 545 85 546
rect 45 540 85 541
rect 45 537 85 538
rect 45 522 85 523
rect 45 519 85 520
rect 45 514 85 515
rect 45 511 85 512
rect 45 478 85 479
rect 282 485 322 486
rect 282 482 322 483
rect 45 475 85 476
rect 282 477 322 478
rect 282 474 322 475
rect 45 460 85 461
rect 45 457 85 458
rect 45 452 85 453
rect 282 459 322 460
rect 282 456 322 457
rect 45 449 85 450
rect 282 451 322 452
rect 282 448 322 449
rect 45 417 85 418
rect 45 414 85 415
rect 45 409 85 410
rect 45 406 85 407
rect 45 262 85 263
rect 45 259 85 260
rect 45 244 85 245
rect 45 241 85 242
rect 45 236 85 237
rect 45 233 85 234
rect 247 231 287 232
rect 247 228 287 229
rect 247 213 287 214
rect 247 210 287 211
rect 247 205 287 206
rect 247 202 287 203
rect 45 194 85 195
rect 45 191 85 192
rect 45 186 85 187
rect 45 183 85 184
rect 46 51 86 52
rect 46 48 86 49
rect 46 43 86 44
rect 46 40 86 41
rect 220 32 260 33
rect 220 29 260 30
rect 220 24 260 25
rect 220 21 260 22
<< ndcontact >>
rect 107 931 207 935
rect 107 923 207 927
rect 107 913 207 917
rect 107 905 207 909
rect 107 897 207 901
rect 107 887 207 891
rect 107 879 207 883
rect 107 871 207 875
rect 107 825 187 829
rect 107 817 187 821
rect 107 809 187 813
rect 389 811 489 815
rect 389 803 489 807
rect 107 799 187 803
rect 107 791 187 795
rect 389 793 489 797
rect 107 783 187 787
rect 389 785 489 789
rect 389 777 489 781
rect 389 767 489 771
rect 107 755 167 759
rect 389 759 489 763
rect 389 751 489 755
rect 107 747 167 751
rect 107 737 167 741
rect 107 729 167 733
rect 107 721 167 725
rect 107 694 147 698
rect 107 686 147 690
rect 107 678 147 682
rect 107 549 187 553
rect 107 541 187 545
rect 107 533 187 537
rect 107 523 187 527
rect 107 515 187 519
rect 107 507 187 511
rect 107 479 167 483
rect 344 486 424 490
rect 107 471 167 475
rect 344 478 424 482
rect 344 470 424 474
rect 107 461 167 465
rect 107 453 167 457
rect 344 460 424 464
rect 107 445 167 449
rect 344 452 424 456
rect 344 444 424 448
rect 107 418 147 422
rect 107 410 147 414
rect 107 402 147 406
rect 107 263 167 267
rect 107 255 167 259
rect 107 245 167 249
rect 107 237 167 241
rect 107 229 167 233
rect 309 232 369 236
rect 309 224 369 228
rect 309 214 369 218
rect 309 206 369 210
rect 107 195 147 199
rect 309 198 369 202
rect 107 187 147 191
rect 107 179 147 183
rect 108 52 148 56
rect 108 44 148 48
rect 108 36 148 40
rect 282 33 322 37
rect 282 25 322 29
rect 282 17 322 21
<< pdcontact >>
rect 45 931 85 935
rect 45 923 85 927
rect 45 913 85 917
rect 45 905 85 909
rect 45 897 85 901
rect 45 887 85 891
rect 45 879 85 883
rect 45 871 85 875
rect 45 825 85 829
rect 45 817 85 821
rect 45 809 85 813
rect 327 811 367 815
rect 327 803 367 807
rect 45 799 85 803
rect 45 791 85 795
rect 327 793 367 797
rect 45 783 85 787
rect 327 785 367 789
rect 327 777 367 781
rect 327 767 367 771
rect 327 759 367 763
rect 45 755 85 759
rect 45 747 85 751
rect 327 751 367 755
rect 45 737 85 741
rect 45 729 85 733
rect 45 721 85 725
rect 45 694 85 698
rect 45 686 85 690
rect 45 678 85 682
rect 45 549 85 553
rect 45 541 85 545
rect 45 533 85 537
rect 45 523 85 527
rect 45 515 85 519
rect 45 507 85 511
rect 282 486 322 490
rect 45 479 85 483
rect 282 478 322 482
rect 45 471 85 475
rect 282 470 322 474
rect 45 461 85 465
rect 282 460 322 464
rect 45 453 85 457
rect 282 452 322 456
rect 45 445 85 449
rect 282 444 322 448
rect 45 418 85 422
rect 45 410 85 414
rect 45 402 85 406
rect 45 263 85 267
rect 45 255 85 259
rect 45 245 85 249
rect 45 237 85 241
rect 45 229 85 233
rect 247 232 287 236
rect 247 224 287 228
rect 247 214 287 218
rect 247 206 287 210
rect 45 195 85 199
rect 247 198 287 202
rect 45 187 85 191
rect 45 179 85 183
rect 46 52 86 56
rect 46 44 86 48
rect 46 36 86 40
rect 220 33 260 37
rect 220 25 260 29
rect 220 17 260 21
<< polysilicon >>
rect 32 928 45 930
rect 85 928 107 930
rect 207 928 210 930
rect 32 910 45 912
rect 85 910 107 912
rect 207 910 210 912
rect 32 902 45 904
rect 85 902 107 904
rect 207 902 210 904
rect 32 884 45 886
rect 85 884 107 886
rect 207 884 210 886
rect 32 876 45 878
rect 85 876 107 878
rect 207 876 210 878
rect 32 822 45 824
rect 85 822 107 824
rect 187 822 190 824
rect 32 814 45 816
rect 85 814 107 816
rect 187 814 190 816
rect 314 808 327 810
rect 367 808 389 810
rect 489 808 492 810
rect 32 796 45 798
rect 85 796 107 798
rect 187 796 190 798
rect 32 788 45 790
rect 85 788 107 790
rect 187 788 190 790
rect 314 790 327 792
rect 367 790 389 792
rect 489 790 492 792
rect 314 782 327 784
rect 367 782 389 784
rect 489 782 492 784
rect 314 764 327 766
rect 367 764 389 766
rect 489 764 492 766
rect 314 756 327 758
rect 367 756 389 758
rect 489 756 492 758
rect 32 752 45 754
rect 85 752 107 754
rect 167 752 170 754
rect 32 734 45 736
rect 85 734 107 736
rect 167 734 170 736
rect 32 726 45 728
rect 85 726 107 728
rect 167 726 170 728
rect 32 691 45 693
rect 85 691 107 693
rect 147 691 150 693
rect 32 683 45 685
rect 85 683 107 685
rect 147 683 150 685
rect 32 546 45 548
rect 85 546 107 548
rect 187 546 190 548
rect 32 538 45 540
rect 85 538 107 540
rect 187 538 190 540
rect 32 520 45 522
rect 85 520 107 522
rect 187 520 190 522
rect 32 512 45 514
rect 85 512 107 514
rect 187 512 190 514
rect 269 483 282 485
rect 322 483 344 485
rect 424 483 427 485
rect 32 476 45 478
rect 85 476 107 478
rect 167 476 170 478
rect 269 475 282 477
rect 322 475 344 477
rect 424 475 427 477
rect 32 458 45 460
rect 85 458 107 460
rect 167 458 170 460
rect 269 457 282 459
rect 322 457 344 459
rect 424 457 427 459
rect 32 450 45 452
rect 85 450 107 452
rect 167 450 170 452
rect 269 449 282 451
rect 322 449 344 451
rect 424 449 427 451
rect 32 415 45 417
rect 85 415 107 417
rect 147 415 150 417
rect 32 407 45 409
rect 85 407 107 409
rect 147 407 150 409
rect 32 260 45 262
rect 85 260 107 262
rect 167 260 170 262
rect 32 242 45 244
rect 85 242 107 244
rect 167 242 170 244
rect 32 234 45 236
rect 85 234 107 236
rect 167 234 170 236
rect 234 229 247 231
rect 287 229 309 231
rect 369 229 372 231
rect 234 211 247 213
rect 287 211 309 213
rect 369 211 372 213
rect 234 203 247 205
rect 287 203 309 205
rect 369 203 372 205
rect 32 192 45 194
rect 85 192 107 194
rect 147 192 150 194
rect 32 184 45 186
rect 85 184 107 186
rect 147 184 150 186
rect 33 49 46 51
rect 86 49 108 51
rect 148 49 151 51
rect 33 41 46 43
rect 86 41 108 43
rect 148 41 151 43
rect 207 30 220 32
rect 260 30 282 32
rect 322 30 325 32
rect 207 22 220 24
rect 260 22 282 24
rect 322 22 325 24
<< polycontact >>
rect 28 927 32 931
rect 28 909 32 913
rect 28 901 32 905
rect 28 883 32 887
rect 28 875 32 879
rect 28 821 32 825
rect 28 813 32 817
rect 310 807 314 811
rect 28 795 32 799
rect 28 787 32 791
rect 310 789 314 793
rect 310 781 314 785
rect 310 763 314 767
rect 28 751 32 755
rect 310 755 314 759
rect 28 733 32 737
rect 28 725 32 729
rect 28 690 32 694
rect 28 682 32 686
rect 28 545 32 549
rect 28 537 32 541
rect 28 519 32 523
rect 28 511 32 515
rect 28 475 32 479
rect 265 482 269 486
rect 265 474 269 478
rect 28 457 32 461
rect 28 449 32 453
rect 265 456 269 460
rect 265 448 269 452
rect 28 414 32 418
rect 28 406 32 410
rect 28 259 32 263
rect 28 241 32 245
rect 28 233 32 237
rect 230 228 234 232
rect 230 210 234 214
rect 230 202 234 206
rect 28 191 32 195
rect 28 183 32 187
rect 29 48 33 52
rect 29 40 33 44
rect 203 29 207 33
rect 203 21 207 25
<< metal1 >>
rect 23 927 28 931
rect 37 927 41 952
rect 85 931 93 935
rect 207 931 218 935
rect 36 923 45 927
rect 23 909 28 913
rect 37 909 41 923
rect 89 917 93 931
rect 85 913 93 917
rect 101 923 107 927
rect 101 917 105 923
rect 101 913 107 917
rect 36 905 45 909
rect 23 901 28 905
rect 23 883 28 887
rect 37 883 41 905
rect 89 901 93 913
rect 85 897 94 901
rect 101 897 107 901
rect 89 891 93 897
rect 85 887 93 891
rect 101 891 105 897
rect 101 887 107 891
rect 36 879 45 883
rect 23 875 28 879
rect 24 821 28 825
rect 37 821 41 879
rect 89 875 93 887
rect 85 871 107 875
rect 97 859 101 871
rect 97 855 304 859
rect 85 825 93 829
rect 187 825 216 829
rect 36 817 45 821
rect 24 813 28 817
rect 23 795 28 799
rect 37 795 41 817
rect 89 813 93 825
rect 85 809 94 813
rect 101 809 107 813
rect 300 811 304 855
rect 89 803 93 809
rect 85 799 93 803
rect 101 803 105 809
rect 300 807 310 811
rect 317 807 321 824
rect 617 816 621 959
rect 593 815 621 816
rect 367 811 375 815
rect 489 811 621 815
rect 300 806 304 807
rect 317 803 327 807
rect 101 799 107 803
rect 36 791 45 795
rect 23 787 28 791
rect 37 759 41 791
rect 89 787 93 799
rect 212 789 310 793
rect 317 789 321 803
rect 371 797 375 811
rect 593 809 621 811
rect 367 793 375 797
rect 383 803 389 807
rect 383 797 387 803
rect 383 793 389 797
rect 85 783 107 787
rect 97 778 101 783
rect 212 778 216 789
rect 317 785 327 789
rect 97 774 216 778
rect 231 781 310 785
rect 36 755 45 759
rect 167 755 216 759
rect 24 751 28 755
rect 23 733 28 737
rect 37 733 41 755
rect 85 747 93 751
rect 89 741 93 747
rect 85 737 93 741
rect 101 747 107 751
rect 101 741 105 747
rect 101 737 107 741
rect 36 729 45 733
rect 23 725 28 729
rect 24 690 28 694
rect 37 690 41 729
rect 89 725 93 737
rect 85 721 107 725
rect 100 716 104 721
rect 231 716 235 781
rect 100 712 235 716
rect 244 763 310 767
rect 317 763 321 785
rect 371 781 375 793
rect 367 777 376 781
rect 383 777 389 781
rect 371 771 375 777
rect 367 767 375 771
rect 383 771 387 777
rect 383 767 389 771
rect 85 694 93 698
rect 147 694 217 698
rect 36 686 45 690
rect 24 682 28 686
rect 37 658 41 686
rect 89 682 93 694
rect 85 678 107 682
rect 100 673 104 678
rect 244 673 248 763
rect 317 759 327 763
rect 306 755 310 759
rect 100 669 248 673
rect 317 658 321 759
rect 371 755 375 767
rect 367 751 389 755
rect 379 709 383 751
rect 379 705 575 709
rect 571 698 575 705
rect 617 685 621 809
rect 536 681 621 685
rect 37 654 321 658
rect 0 545 28 549
rect 37 545 41 654
rect 85 549 93 553
rect 187 549 207 553
rect 36 541 45 545
rect 6 537 28 541
rect 14 519 28 523
rect 37 519 41 541
rect 89 537 93 549
rect 85 533 94 537
rect 101 533 107 537
rect 89 527 93 533
rect 85 523 93 527
rect 101 527 105 533
rect 101 523 107 527
rect 36 515 45 519
rect 22 511 28 515
rect 37 483 41 515
rect 89 511 93 523
rect 85 507 107 511
rect 97 494 101 507
rect 97 490 199 494
rect 195 486 199 490
rect 36 479 45 483
rect 167 479 182 483
rect 6 475 28 479
rect 14 457 28 461
rect 37 457 41 479
rect 187 479 188 483
rect 195 482 265 486
rect 273 482 277 496
rect 617 490 621 681
rect 322 486 330 490
rect 424 486 621 490
rect 273 478 282 482
rect 85 471 93 475
rect 89 465 93 471
rect 85 461 93 465
rect 101 471 107 475
rect 192 474 265 478
rect 101 465 105 471
rect 101 461 107 465
rect 36 453 45 457
rect 21 449 28 453
rect 14 414 28 418
rect 37 414 41 453
rect 89 449 93 461
rect 85 445 107 449
rect 99 441 103 445
rect 192 441 196 474
rect 99 437 196 441
rect 206 456 265 460
rect 273 456 277 478
rect 326 474 330 486
rect 322 470 331 474
rect 338 470 344 474
rect 326 464 330 470
rect 322 460 330 464
rect 338 464 342 470
rect 338 460 344 464
rect 85 418 93 422
rect 147 419 183 422
rect 188 419 193 422
rect 147 418 193 419
rect 36 410 45 414
rect 22 406 28 410
rect 37 377 41 410
rect 89 406 93 418
rect 85 402 107 406
rect 96 398 100 402
rect 206 398 210 456
rect 273 452 282 456
rect 259 448 265 452
rect 96 394 210 398
rect 273 377 277 452
rect 326 448 330 460
rect 322 444 344 448
rect 331 396 335 444
rect 617 423 621 486
rect 457 419 621 423
rect 331 392 532 396
rect 37 373 277 377
rect 37 267 41 373
rect 617 341 621 419
rect 444 337 621 341
rect 444 281 448 337
rect 412 277 448 281
rect 36 263 45 267
rect 167 263 185 267
rect 6 259 28 263
rect 14 241 28 245
rect 37 241 41 263
rect 85 255 93 259
rect 89 249 93 255
rect 85 245 93 249
rect 101 255 107 259
rect 101 249 105 255
rect 101 245 107 249
rect 36 237 45 241
rect 22 233 28 237
rect 11 191 28 195
rect 37 191 41 237
rect 89 233 93 245
rect 237 236 241 248
rect 444 236 448 277
rect 85 229 107 233
rect 237 232 247 236
rect 369 232 448 236
rect 97 221 101 229
rect 193 228 230 232
rect 193 221 197 228
rect 97 217 197 221
rect 205 210 230 214
rect 237 210 241 232
rect 287 224 295 228
rect 291 218 295 224
rect 287 214 295 218
rect 303 224 309 228
rect 303 218 307 224
rect 303 214 309 218
rect 85 195 93 199
rect 147 195 185 199
rect 36 187 45 191
rect 6 183 28 187
rect 37 158 41 187
rect 89 183 93 195
rect 85 179 107 183
rect 98 174 102 179
rect 205 174 209 210
rect 237 206 247 210
rect 224 202 230 206
rect 98 170 209 174
rect 237 158 241 206
rect 291 202 295 214
rect 287 198 309 202
rect 299 176 303 198
rect 299 172 411 176
rect 37 154 241 158
rect 6 48 29 52
rect 37 48 41 154
rect 444 56 448 232
rect 86 52 94 56
rect 148 52 448 56
rect 37 44 46 48
rect 23 40 29 44
rect 37 -7 41 44
rect 90 40 94 52
rect 86 36 108 40
rect 326 37 330 52
rect 99 33 103 36
rect 260 33 268 37
rect 322 33 330 37
rect 99 29 203 33
rect 211 25 220 29
rect 197 21 203 25
rect 264 21 268 33
rect 260 17 282 21
rect 271 4 275 17
rect 271 0 389 4
<< m2contact >>
rect 218 931 223 936
rect 216 825 221 830
rect 216 755 221 760
rect 217 694 222 699
rect 531 681 536 686
rect 207 548 212 553
rect 182 478 187 483
rect 183 419 188 424
rect 452 419 457 424
rect 407 277 412 282
rect 185 263 190 268
rect 185 195 190 200
<< metal2 >>
rect 218 936 221 947
rect 218 836 221 931
rect 217 830 221 836
rect 217 760 221 825
rect 217 699 221 755
rect 217 685 221 694
rect 217 681 531 685
rect 207 499 211 548
rect 183 495 211 499
rect 183 483 187 495
rect 183 424 187 478
rect 188 419 452 423
rect 185 277 407 281
rect 185 268 189 277
rect 185 200 189 263
<< labels >>
rlabel metal1 197 21 200 25 1 g1
rlabel metal1 225 202 228 206 1 g2
rlabel metal1 260 448 263 452 1 g3
rlabel metal1 306 755 309 759 1 g4
rlabel metal1 24 40 27 44 1 g0
rlabel metal1 23 875 26 879 1 g0
rlabel metal1 23 787 26 791 1 g1
rlabel metal1 23 725 26 729 1 g2
rlabel metal1 24 682 27 686 1 g3
rlabel metal1 23 511 26 515 1 g0
rlabel metal1 24 449 27 453 1 g1
rlabel metal1 24 406 27 410 1 g2
rlabel metal1 24 183 27 187 1 g1
rlabel metal1 24 48 27 52 1 p1
rlabel metal1 24 191 27 195 1 p2
rlabel metal1 24 414 27 418 1 p3
rlabel metal1 24 457 27 461 1 p2
rlabel metal1 24 475 27 479 1 p3
rlabel metal1 23 519 26 523 1 p1
rlabel metal1 23 537 26 541 1 p2
rlabel metal1 23 545 26 549 1 p3
rlabel metal1 24 690 27 694 1 p4
rlabel metal1 23 733 26 737 1 p3
rlabel metal1 24 751 27 755 1 p4
rlabel metal1 23 795 26 799 1 p2
rlabel metal1 24 813 27 817 1 p3
rlabel metal1 24 821 27 825 1 p4
rlabel metal1 384 0 388 4 1 c2
rlabel metal1 405 172 409 176 1 c3
rlabel metal1 518 392 522 396 1 c4
rlabel metal1 562 705 566 709 1 c5
rlabel metal1 23 901 26 905 1 p2
rlabel metal1 23 883 26 887 1 p1
rlabel metal1 23 909 26 913 1 p3
rlabel metal1 23 927 26 931 1 p4
rlabel metal1 24 233 27 237 1 g0
rlabel metal1 24 241 27 245 1 p1
rlabel metal1 23 259 26 263 1 p2
rlabel metal1 37 -7 41 -3 1 vdd
rlabel metal1 617 955 621 959 6 gnd
<< end >>
