magic
tech scmos
timestamp 1763524194
<< nwell >>
rect 264 235 288 291
rect 384 234 408 290
rect 311 130 359 222
rect 86 -26 110 30
rect 206 -27 230 29
rect 133 -131 181 -39
<< ntransistor >>
rect 275 299 277 319
rect 395 298 397 318
rect 322 74 324 114
rect 330 74 332 114
rect 338 74 340 114
rect 346 74 348 114
rect 97 38 99 58
rect 217 37 219 57
rect 144 -187 146 -147
rect 152 -187 154 -147
rect 160 -187 162 -147
rect 168 -187 170 -147
<< ptransistor >>
rect 275 245 277 285
rect 395 244 397 284
rect 322 136 324 216
rect 330 136 332 216
rect 338 136 340 216
rect 346 136 348 216
rect 97 -16 99 24
rect 217 -17 219 23
rect 144 -125 146 -45
rect 152 -125 154 -45
rect 160 -125 162 -45
rect 168 -125 170 -45
<< ndiffusion >>
rect 274 299 275 319
rect 277 299 278 319
rect 394 298 395 318
rect 397 298 398 318
rect 321 74 322 114
rect 324 74 325 114
rect 329 74 330 114
rect 332 74 333 114
rect 337 74 338 114
rect 340 74 341 114
rect 345 74 346 114
rect 348 74 349 114
rect 96 38 97 58
rect 99 38 100 58
rect 216 37 217 57
rect 219 37 220 57
rect 143 -187 144 -147
rect 146 -187 147 -147
rect 151 -187 152 -147
rect 154 -187 155 -147
rect 159 -187 160 -147
rect 162 -187 163 -147
rect 167 -187 168 -147
rect 170 -187 171 -147
<< pdiffusion >>
rect 274 245 275 285
rect 277 245 278 285
rect 394 244 395 284
rect 397 244 398 284
rect 321 136 322 216
rect 324 136 325 216
rect 329 136 330 216
rect 332 136 333 216
rect 337 136 338 216
rect 340 136 341 216
rect 345 136 346 216
rect 348 136 349 216
rect 96 -16 97 24
rect 99 -16 100 24
rect 216 -17 217 23
rect 219 -17 220 23
rect 143 -125 144 -45
rect 146 -125 147 -45
rect 151 -125 152 -45
rect 154 -125 155 -45
rect 159 -125 160 -45
rect 162 -125 163 -45
rect 167 -125 168 -45
rect 170 -125 171 -45
<< ndcontact >>
rect 270 299 274 319
rect 278 299 282 319
rect 390 298 394 318
rect 398 298 402 318
rect 317 74 321 114
rect 325 74 329 114
rect 333 74 337 114
rect 341 74 345 114
rect 349 74 353 114
rect 92 38 96 58
rect 100 38 104 58
rect 212 37 216 57
rect 220 37 224 57
rect 139 -187 143 -147
rect 147 -187 151 -147
rect 155 -187 159 -147
rect 163 -187 167 -147
rect 171 -187 175 -147
<< pdcontact >>
rect 270 245 274 285
rect 278 245 282 285
rect 390 244 394 284
rect 398 244 402 284
rect 317 136 321 216
rect 325 136 329 216
rect 333 136 337 216
rect 341 136 345 216
rect 349 136 353 216
rect 92 -16 96 24
rect 100 -16 104 24
rect 212 -17 216 23
rect 220 -17 224 23
rect 139 -125 143 -45
rect 147 -125 151 -45
rect 155 -125 159 -45
rect 163 -125 167 -45
rect 171 -125 175 -45
<< polysilicon >>
rect 275 319 277 322
rect 395 318 397 321
rect 275 285 277 299
rect 395 284 397 298
rect 275 242 277 245
rect 395 241 397 244
rect 322 216 324 229
rect 330 216 332 229
rect 338 216 340 229
rect 346 216 348 229
rect 322 133 324 136
rect 330 125 332 136
rect 322 123 332 125
rect 338 125 340 136
rect 346 133 348 136
rect 338 123 348 125
rect 322 114 324 123
rect 330 114 332 117
rect 338 114 340 117
rect 346 114 348 123
rect 322 71 324 74
rect 330 66 332 74
rect 324 64 332 66
rect 338 66 340 74
rect 346 71 348 74
rect 338 64 347 66
rect 97 58 99 61
rect 217 57 219 60
rect 97 24 99 38
rect 217 23 219 37
rect 97 -19 99 -16
rect 217 -20 219 -17
rect 144 -45 146 -32
rect 152 -45 154 -32
rect 160 -45 162 -32
rect 168 -45 170 -32
rect 144 -128 146 -125
rect 152 -136 154 -125
rect 144 -138 154 -136
rect 160 -136 162 -125
rect 168 -128 170 -125
rect 160 -138 170 -136
rect 144 -147 146 -138
rect 152 -147 154 -144
rect 160 -147 162 -144
rect 168 -147 170 -138
rect 144 -190 146 -187
rect 152 -195 154 -187
rect 146 -197 154 -195
rect 160 -195 162 -187
rect 168 -190 170 -187
rect 160 -197 169 -195
<< polycontact >>
rect 277 292 281 296
rect 397 291 401 295
rect 321 229 325 233
rect 329 229 333 233
rect 337 229 341 233
rect 345 229 349 233
rect 320 63 324 67
rect 347 63 351 67
rect 99 31 103 35
rect 219 30 223 34
rect 143 -32 147 -28
rect 151 -32 155 -28
rect 159 -32 163 -28
rect 167 -32 171 -28
rect 142 -198 146 -194
rect 169 -198 173 -194
<< metal1 >>
rect 247 323 283 327
rect 247 219 251 323
rect 278 319 282 323
rect 270 296 274 299
rect 337 296 341 352
rect 398 323 402 324
rect 398 319 424 323
rect 398 318 402 319
rect 256 292 274 296
rect 281 292 341 296
rect 390 295 394 298
rect 257 230 261 292
rect 270 285 274 292
rect 307 261 333 265
rect 278 239 282 245
rect 291 239 296 240
rect 264 235 296 239
rect 307 230 311 261
rect 322 235 325 249
rect 257 226 311 230
rect 321 233 325 235
rect 329 233 333 261
rect 337 233 341 292
rect 345 291 394 295
rect 401 291 412 295
rect 345 233 349 291
rect 362 286 366 291
rect 390 284 394 291
rect 370 225 374 239
rect 398 238 402 244
rect 420 239 424 319
rect 434 251 438 333
rect 433 247 484 251
rect 384 234 411 238
rect 407 225 411 234
rect 434 225 438 247
rect 333 221 438 225
rect 247 215 294 219
rect 333 216 337 221
rect 317 123 321 136
rect 349 123 353 136
rect 159 119 353 123
rect 69 62 105 66
rect 69 -42 73 62
rect 100 58 104 62
rect 92 35 96 38
rect 159 35 163 119
rect 317 114 321 119
rect 349 114 353 119
rect 220 62 224 63
rect 220 58 246 62
rect 220 57 224 58
rect 78 31 96 35
rect 103 31 163 35
rect 212 34 216 37
rect 79 -31 83 31
rect 92 24 96 31
rect 129 0 155 4
rect 100 -22 104 -16
rect 113 -22 118 -21
rect 86 -26 118 -22
rect 129 -31 133 0
rect 144 -26 147 -12
rect 79 -35 133 -31
rect 143 -28 147 -26
rect 151 -28 155 0
rect 159 -28 163 31
rect 167 30 216 34
rect 223 30 234 34
rect 167 -28 171 30
rect 184 25 188 30
rect 212 23 216 30
rect 192 -36 196 -22
rect 220 -23 224 -17
rect 242 -22 246 58
rect 256 -10 260 72
rect 333 63 337 74
rect 321 40 324 63
rect 347 59 350 63
rect 362 40 365 158
rect 321 37 365 40
rect 480 -10 484 247
rect 255 -14 484 -10
rect 206 -27 233 -23
rect 229 -36 233 -27
rect 256 -36 260 -14
rect 155 -40 260 -36
rect 69 -46 116 -42
rect 155 -45 159 -40
rect 139 -138 143 -125
rect 171 -138 175 -125
rect 101 -142 175 -138
rect 139 -147 143 -142
rect 171 -147 175 -142
rect 155 -198 159 -187
rect 143 -221 146 -198
rect 169 -202 172 -198
rect 184 -221 187 -103
rect 143 -224 187 -221
<< m2contact >>
rect 291 240 297 246
rect 321 249 326 254
rect 362 280 368 286
rect 370 239 376 245
rect 419 233 425 239
rect 294 214 300 220
rect 362 158 367 163
rect 113 -21 119 -15
rect 143 -12 148 -7
rect 184 19 190 25
rect 192 -22 198 -16
rect 332 57 338 63
rect 347 54 352 59
rect 241 -28 247 -22
rect 116 -47 122 -41
rect 184 -103 189 -98
rect 154 -204 160 -198
rect 169 -207 174 -202
<< metal2 >>
rect 412 342 415 350
rect 322 339 415 342
rect 322 254 325 339
rect 363 257 366 280
rect 297 240 370 244
rect 412 214 415 339
rect 234 81 237 89
rect 144 78 237 81
rect 144 -7 147 78
rect 185 -4 188 19
rect 119 -21 192 -17
rect 234 -47 237 78
rect 294 36 298 214
rect 382 211 415 214
rect 363 163 366 171
rect 333 36 337 57
rect 348 49 351 54
rect 382 49 385 211
rect 421 203 425 233
rect 348 46 385 49
rect 390 199 425 203
rect 294 35 339 36
rect 390 35 394 199
rect 294 32 394 35
rect 333 31 394 32
rect 116 -225 120 -47
rect 204 -50 237 -47
rect 185 -98 188 -90
rect 155 -225 159 -204
rect 170 -212 173 -207
rect 204 -212 207 -50
rect 243 -58 247 -28
rect 170 -215 207 -212
rect 212 -62 247 -58
rect 212 -135 216 -62
rect 389 -135 393 31
rect 212 -139 393 -135
rect 116 -226 161 -225
rect 212 -226 216 -139
rect 116 -229 216 -226
rect 155 -230 216 -229
rect 211 -236 215 -230
<< m3contact >>
rect 362 252 367 257
rect 184 -9 189 -4
rect 361 171 367 178
rect 183 -90 189 -83
<< metal3 >>
rect 363 178 366 252
rect 185 -83 188 -9
<< labels >>
rlabel metal1 337 346 341 351 1 a
rlabel metal1 434 328 438 333 7 vdd
rlabel metal2 389 24 393 28 1 gnd
rlabel metal2 412 346 415 350 5 b
rlabel metal1 308 119 311 123 1 axorb
rlabel metal2 234 83 237 89 1 c
rlabel metal1 101 -142 104 -138 1 axorbxorc
<< end >>
