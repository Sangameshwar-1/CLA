* Comprehensive Test Bench for 5-bit Carry Lookahead Adder (CMOS-static-2)
* Tests multiple addition cases with detailed verification

.include "TSMC_180nm.txt"

* Technology parameters (CMOS-static-2)
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_P=0.18u
.param width_N=0.09u

* Include all subcircuit files (order matters!)
.include "inv.cir"
.include "nand_2.cir"
.include "nand_3.cir"
.include "nand_4.cir"
.include "nand_5.cir"
.include "xor.cir"
.include "gi_bar.cir"
.include "pi.cir"
.include "si.cir"
.include "carry.cir"

* Power supplies
Vdd vdd 0 DC {SUPPLY}

* ============================================
* TEST 1: 0+0=0 (00000+00000=00000)
* ============================================
Va0_t1 a0_t1 0 DC 0
Va1_t1 a1_t1 0 DC 0
Va2_t1 a2_t1 0 DC 0
Va3_t1 a3_t1 0 DC 0
Va4_t1 a4_t1 0 DC 0
Vb0_t1 b0_t1 0 DC 0
Vb1_t1 b1_t1 0 DC 0
Vb2_t1 b2_t1 0 DC 0
Vb3_t1 b3_t1 0 DC 0
Vb4_t1 b4_t1 0 DC 0

* Use 'gi' as subcircuit name (not 'gi_bar')
Xgi_bar_t1 a0_t1 a1_t1 a2_t1 a3_t1 a4_t1 b0_t1 b1_t1 b2_t1 b3_t1 b4_t1 g0bar_t1 g1bar_t1 g2bar_t1 g3bar_t1 g4bar_t1 vdd 0 gi
Xpi_t1 a0_t1 a1_t1 a2_t1 a3_t1 a4_t1 b0_t1 b1_t1 b2_t1 b3_t1 b4_t1 p0_t1 p1_t1 p2_t1 p3_t1 p4_t1 vdd 0 pi
Xcarry_t1 p0_t1 p1_t1 p2_t1 p3_t1 p4_t1 g0bar_t1 g1bar_t1 g2bar_t1 g3bar_t1 g4bar_t1 c1_t1 c2_t1 c3_t1 c4_t1 c5_t1 vdd 0 carry
Vc0_t1 c0_t1 0 DC 0
Xsi_t1 p0_t1 p1_t1 p2_t1 p3_t1 p4_t1 c0_t1 c1_t1 c2_t1 c3_t1 c4_t1 s0_t1 s1_t1 s2_t1 s3_t1 s4_t1 vdd 0 si

* ============================================
* TEST 2: 1+1=2 (00001+00001=00010)
* ============================================
Va0_t2 a0_t2 0 DC {SUPPLY}
Va1_t2 a1_t2 0 DC 0
Va2_t2 a2_t2 0 DC 0
Va3_t2 a3_t2 0 DC 0
Va4_t2 a4_t2 0 DC 0
Vb0_t2 b0_t2 0 DC {SUPPLY}
Vb1_t2 b1_t2 0 DC 0
Vb2_t2 b2_t2 0 DC 0
Vb3_t2 b3_t2 0 DC 0
Vb4_t2 b4_t2 0 DC 0

Xgi_bar_t2 a0_t2 a1_t2 a2_t2 a3_t2 a4_t2 b0_t2 b1_t2 b2_t2 b3_t2 b4_t2 g0bar_t2 g1bar_t2 g2bar_t2 g3bar_t2 g4bar_t2 vdd 0 gi
Xpi_t2 a0_t2 a1_t2 a2_t2 a3_t2 a4_t2 b0_t2 b1_t2 b2_t2 b3_t2 b4_t2 p0_t2 p1_t2 p2_t2 p3_t2 p4_t2 vdd 0 pi
Xcarry_t2 p0_t2 p1_t2 p2_t2 p3_t2 p4_t2 g0bar_t2 g1bar_t2 g2bar_t2 g3bar_t2 g4bar_t2 c1_t2 c2_t2 c3_t2 c4_t2 c5_t2 vdd 0 carry
Vc0_t2 c0_t2 0 DC 0
Xsi_t2 p0_t2 p1_t2 p2_t2 p3_t2 p4_t2 c0_t2 c1_t2 c2_t2 c3_t2 c4_t2 s0_t2 s1_t2 s2_t2 s3_t2 s4_t2 vdd 0 si

* ============================================
* TEST 3: 7+8=15 (00111+01000=01111)
* ============================================
Va0_t3 a0_t3 0 DC {SUPPLY}
Va1_t3 a1_t3 0 DC {SUPPLY}
Va2_t3 a2_t3 0 DC {SUPPLY}
Va3_t3 a3_t3 0 DC 0
Va4_t3 a4_t3 0 DC 0
Vb0_t3 b0_t3 0 DC 0
Vb1_t3 b1_t3 0 DC 0
Vb2_t3 b2_t3 0 DC 0
Vb3_t3 b3_t3 0 DC {SUPPLY}
Vb4_t3 b4_t3 0 DC 0

Xgi_bar_t3 a0_t3 a1_t3 a2_t3 a3_t3 a4_t3 b0_t3 b1_t3 b2_t3 b3_t3 b4_t3 g0bar_t3 g1bar_t3 g2bar_t3 g3bar_t3 g4bar_t3 vdd 0 gi
Xpi_t3 a0_t3 a1_t3 a2_t3 a3_t3 a4_t3 b0_t3 b1_t3 b2_t3 b3_t3 b4_t3 p0_t3 p1_t3 p2_t3 p3_t3 p4_t3 vdd 0 pi
Xcarry_t3 p0_t3 p1_t3 p2_t3 p3_t3 p4_t3 g0bar_t3 g1bar_t3 g2bar_t3 g3bar_t3 g4bar_t3 c1_t3 c2_t3 c3_t3 c4_t3 c5_t3 vdd 0 carry
Vc0_t3 c0_t3 0 DC 0
Xsi_t3 p0_t3 p1_t3 p2_t3 p3_t3 p4_t3 c0_t3 c1_t3 c2_t3 c3_t3 c4_t3 s0_t3 s1_t3 s2_t3 s3_t3 s4_t3 vdd 0 si

* ============================================
* TEST 4: 15+1=16 (01111+00001=10000)
* ============================================
Va0_t4 a0_t4 0 DC {SUPPLY}
Va1_t4 a1_t4 0 DC {SUPPLY}
Va2_t4 a2_t4 0 DC {SUPPLY}
Va3_t4 a3_t4 0 DC {SUPPLY}
Va4_t4 a4_t4 0 DC 0
Vb0_t4 b0_t4 0 DC {SUPPLY}
Vb1_t4 b1_t4 0 DC 0
Vb2_t4 b2_t4 0 DC 0
Vb3_t4 b3_t4 0 DC 0
Vb4_t4 b4_t4 0 DC 0

Xgi_bar_t4 a0_t4 a1_t4 a2_t4 a3_t4 a4_t4 b0_t4 b1_t4 b2_t4 b3_t4 b4_t4 g0bar_t4 g1bar_t4 g2bar_t4 g3bar_t4 g4bar_t4 vdd 0 gi
Xpi_t4 a0_t4 a1_t4 a2_t4 a3_t4 a4_t4 b0_t4 b1_t4 b2_t4 b3_t4 b4_t4 p0_t4 p1_t4 p2_t4 p3_t4 p4_t4 vdd 0 pi
Xcarry_t4 p0_t4 p1_t4 p2_t4 p3_t4 p4_t4 g0bar_t4 g1bar_t4 g2bar_t4 g3bar_t4 g4bar_t4 c1_t4 c2_t4 c3_t4 c4_t4 c5_t4 vdd 0 carry
Vc0_t4 c0_t4 0 DC 0
Xsi_t4 p0_t4 p1_t4 p2_t4 p3_t4 p4_t4 c0_t4 c1_t4 c2_t4 c3_t4 c4_t4 s0_t4 s1_t4 s2_t4 s3_t4 s4_t4 vdd 0 si

* ============================================
* TEST 5: 31+31=62 (11111+11111=11110, Cout=1)
* ============================================
Va0_t5 a0_t5 0 DC {SUPPLY}
Va1_t5 a1_t5 0 DC {SUPPLY}
Va2_t5 a2_t5 0 DC {SUPPLY}
Va3_t5 a3_t5 0 DC {SUPPLY}
Va4_t5 a4_t5 0 DC {SUPPLY}
Vb0_t5 b0_t5 0 DC {SUPPLY}
Vb1_t5 b1_t5 0 DC {SUPPLY}
Vb2_t5 b2_t5 0 DC {SUPPLY}
Vb3_t5 b3_t5 0 DC {SUPPLY}
Vb4_t5 b4_t5 0 DC {SUPPLY}

Xgi_bar_t5 a0_t5 a1_t5 a2_t5 a3_t5 a4_t5 b0_t5 b1_t5 b2_t5 b3_t5 b4_t5 g0bar_t5 g1bar_t5 g2bar_t5 g3bar_t5 g4bar_t5 vdd 0 gi
Xpi_t5 a0_t5 a1_t5 a2_t5 a3_t5 a4_t5 b0_t5 b1_t5 b2_t5 b3_t5 b4_t5 p0_t5 p1_t5 p2_t5 p3_t5 p4_t5 vdd 0 pi
Xcarry_t5 p0_t5 p1_t5 p2_t5 p3_t5 p4_t5 g0bar_t5 g1bar_t5 g2bar_t5 g3bar_t5 g4bar_t5 c1_t5 c2_t5 c3_t5 c4_t5 c5_t5 vdd 0 carry
Vc0_t5 c0_t5 0 DC 0
Xsi_t5 p0_t5 p1_t5 p2_t5 p3_t5 p4_t5 c0_t5 c1_t5 c2_t5 c3_t5 c4_t5 s0_t5 s1_t5 s2_t5 s3_t5 s4_t5 vdd 0 si

* ============================================
* TEST 6: 10+5=15 (01010+00101=01111)
* ============================================
Va0_t6 a0_t6 0 DC 0
Va1_t6 a1_t6 0 DC {SUPPLY}
Va2_t6 a2_t6 0 DC 0
Va3_t6 a3_t6 0 DC {SUPPLY}
Va4_t6 a4_t6 0 DC 0
Vb0_t6 b0_t6 0 DC {SUPPLY}
Vb1_t6 b1_t6 0 DC 0
Vb2_t6 b2_t6 0 DC {SUPPLY}
Vb3_t6 b3_t6 0 DC 0
Vb4_t6 b4_t6 0 DC 0

Xgi_bar_t6 a0_t6 a1_t6 a2_t6 a3_t6 a4_t6 b0_t6 b1_t6 b2_t6 b3_t6 b4_t6 g0bar_t6 g1bar_t6 g2bar_t6 g3bar_t6 g4bar_t6 vdd 0 gi
Xpi_t6 a0_t6 a1_t6 a2_t6 a3_t6 a4_t6 b0_t6 b1_t6 b2_t6 b3_t6 b4_t6 p0_t6 p1_t6 p2_t6 p3_t6 p4_t6 vdd 0 pi
Xcarry_t6 p0_t6 p1_t6 p2_t6 p3_t6 p4_t6 g0bar_t6 g1bar_t6 g2bar_t6 g3bar_t6 g4bar_t6 c1_t6 c2_t6 c3_t6 c4_t6 c5_t6 vdd 0 carry
Vc0_t6 c0_t6 0 DC 0
Xsi_t6 p0_t6 p1_t6 p2_t6 p3_t6 p4_t6 c0_t6 c1_t6 c2_t6 c3_t6 c4_t6 s0_t6 s1_t6 s2_t6 s3_t6 s4_t6 vdd 0 si

* ============================================
* TEST 7: 16+16=32 (10000+10000=00000, Cout=1)
* ============================================
Va0_t7 a0_t7 0 DC 0
Va1_t7 a1_t7 0 DC 0
Va2_t7 a2_t7 0 DC 0
Va3_t7 a3_t7 0 DC 0
Va4_t7 a4_t7 0 DC {SUPPLY}
Vb0_t7 b0_t7 0 DC 0
Vb1_t7 b1_t7 0 DC 0
Vb2_t7 b2_t7 0 DC 0
Vb3_t7 b3_t7 0 DC 0
Vb4_t7 b4_t7 0 DC {SUPPLY}

Xgi_bar_t7 a0_t7 a1_t7 a2_t7 a3_t7 a4_t7 b0_t7 b1_t7 b2_t7 b3_t7 b4_t7 g0bar_t7 g1bar_t7 g2bar_t7 g3bar_t7 g4bar_t7 vdd 0 gi
Xpi_t7 a0_t7 a1_t7 a2_t7 a3_t7 a4_t7 b0_t7 b1_t7 b2_t7 b3_t7 b4_t7 p0_t7 p1_t7 p2_t7 p3_t7 p4_t7 vdd 0 pi
Xcarry_t7 p0_t7 p1_t7 p2_t7 p3_t7 p4_t7 g0bar_t7 g1bar_t7 g2bar_t7 g3bar_t7 g4bar_t7 c1_t7 c2_t7 c3_t7 c4_t7 c5_t7 vdd 0 carry
Vc0_t7 c0_t7 0 DC 0
Xsi_t7 p0_t7 p1_t7 p2_t7 p3_t7 p4_t7 c0_t7 c1_t7 c2_t7 c3_t7 c4_t7 s0_t7 s1_t7 s2_t7 s3_t7 s4_t7 vdd 0 si

* Simulation options
.options METHOD=GEAR MAXORD=2
.options ABSTOL=1e-8 RELTOL=1e-4 VNTOL=1e-5
.options ITL1=500 ITL2=200 ITL4=100
.options TEMP=27

* DC operating point analysis
.op

* Control block
.control
set hcopydevtype=postscript
option numdgt=7

op

echo ""
echo "================================================================"
echo "  5-BIT CARRY LOOKAHEAD ADDER TEST SUITE"
echo "  TSMC 180nm Process (CMOS-static-2)"
echo "================================================================"
echo ""

* Test results display
echo "TEST 1: 0+0=0 (00000+00000=00000)"
echo "Expected: S=00000, Cout=0"
echo "----------------------------------------------------------------"
print v(a4_t1) v(a3_t1) v(a2_t1) v(a1_t1) v(a0_t1)
print v(b4_t1) v(b3_t1) v(b2_t1) v(b1_t1) v(b0_t1)
print v(s4_t1) v(s3_t1) v(s2_t1) v(s1_t1) v(s0_t1) v(c5_t1)
echo ""

echo "TEST 2: 1+1=2 (00001+00001=00010)"
echo "Expected: S=00010, Cout=0"
echo "----------------------------------------------------------------"
print v(a4_t2) v(a3_t2) v(a2_t2) v(a1_t2) v(a0_t2)
print v(b4_t2) v(b3_t2) v(b2_t2) v(b1_t2) v(b0_t2)
print v(s4_t2) v(s3_t2) v(s2_t2) v(s1_t2) v(s0_t2) v(c5_t2)
echo "Carries: C[4:1] ="
print v(c4_t2) v(c3_t2) v(c2_t2) v(c1_t2)
echo ""

echo "TEST 3: 7+8=15 (00111+01000=01111)"
echo "Expected: S=01111, Cout=0"
echo "----------------------------------------------------------------"
print v(a4_t3) v(a3_t3) v(a2_t3) v(a1_t3) v(a0_t3)
print v(b4_t3) v(b3_t3) v(b2_t3) v(b1_t3) v(b0_t3)
print v(s4_t3) v(s3_t3) v(s2_t3) v(s1_t3) v(s0_t3) v(c5_t3)
echo "Carries: C[4:1] ="
print v(c4_t3) v(c3_t3) v(c2_t3) v(c1_t3)
echo ""

echo "TEST 4: 15+1=16 (01111+00001=10000)"
echo "Expected: S=10000, Cout=0"
echo "----------------------------------------------------------------"
print v(a4_t4) v(a3_t4) v(a2_t4) v(a1_t4) v(a0_t4)
print v(b4_t4) v(b3_t4) v(b2_t4) v(b1_t4) v(b0_t4)
print v(s4_t4) v(s3_t4) v(s2_t4) v(s1_t4) v(s0_t4) v(c5_t4)
echo "Carries: C[4:1] ="
print v(c4_t4) v(c3_t4) v(c2_t4) v(c1_t4)
echo ""

echo "TEST 5: 31+31=62 (11111+11111=11110, overflow)"
echo "Expected: S=11110, Cout=1"
echo "----------------------------------------------------------------"
print v(a4_t5) v(a3_t5) v(a2_t5) v(a1_t5) v(a0_t5)
print v(b4_t5) v(b3_t5) v(b2_t5) v(b1_t5) v(b0_t5)
print v(s4_t5) v(s3_t5) v(s2_t5) v(s1_t5) v(s0_t5) v(c5_t5)
echo "Carries: C[4:1] ="
print v(c4_t5) v(c3_t5) v(c2_t5) v(c1_t5)
echo ""

echo "TEST 6: 10+5=15 (01010+00101=01111)"
echo "Expected: S=01111, Cout=0"
echo "----------------------------------------------------------------"
print v(a4_t6) v(a3_t6) v(a2_t6) v(a1_t6) v(a0_t6)
print v(b4_t6) v(b3_t6) v(b2_t6) v(b1_t6) v(b0_t6)
print v(s4_t6) v(s3_t6) v(s2_t6) v(s1_t6) v(s0_t6) v(c5_t6)
echo "Carries: C[4:1] ="
print v(c4_t6) v(c3_t6) v(c2_t6) v(c1_t6)
echo ""

echo "TEST 7: 16+16=32 (10000+10000=00000, overflow)"
echo "Expected: S=00000, Cout=1"
echo "----------------------------------------------------------------"
print v(a4_t7) v(a3_t7) v(a2_t7) v(a1_t7) v(a0_t7)
print v(b4_t7) v(b3_t7) v(b2_t7) v(b1_t7) v(b0_t7)
print v(s4_t7) v(s3_t7) v(s2_t7) v(s1_t7) v(s0_t7) v(c5_t7)
echo "Carries: C[4:1] ="
print v(c4_t7) v(c3_t7) v(c2_t7) v(c1_t7)
echo ""

* Save results
set wr_vecnames
set wr_singlescale
wrdata test_5bit_cla_results.txt v(s4_t1) v(s3_t1) v(s2_t1) v(s1_t1) v(s0_t1) v(c5_t1) v(s4_t2) v(s3_t2) v(s2_t2) v(s1_t2) v(s0_t2) v(c5_t2) v(s4_t5) v(s3_t5) v(s2_t5) v(s1_t5) v(s0_t5) v(c5_t5)

echo "================================================================"
echo "Simulation Complete!"
echo "Results saved to: test_5bit_cla_results.txt"
echo "================================================================"

.endc
.end