magic
tech scmos
timestamp 1763548257
<< nwell >>
rect -18 703 34 735
rect 74 701 126 703
rect -93 665 -41 697
rect 73 669 126 701
rect -21 631 31 663
rect -21 547 31 579
rect 71 545 123 547
rect -96 509 -44 541
rect 70 513 123 545
rect -24 475 28 507
rect -25 392 27 424
rect 67 390 119 392
rect -100 354 -48 386
rect 66 358 119 390
rect -28 320 24 352
rect -28 234 24 266
rect 64 232 116 234
rect -103 196 -51 228
rect 63 200 116 232
rect -31 162 21 194
rect -31 30 21 62
rect 61 28 113 30
rect -106 -8 -54 24
rect 60 -4 113 28
rect -34 -42 18 -10
<< ntransistor >>
rect 50 722 90 724
rect 50 714 90 716
rect 142 690 182 692
rect -25 684 15 686
rect 142 682 182 684
rect -25 676 15 678
rect 47 650 87 652
rect 47 642 87 644
rect 47 566 87 568
rect 47 558 87 560
rect 139 534 179 536
rect -28 528 12 530
rect 139 526 179 528
rect -28 520 12 522
rect 44 494 84 496
rect 44 486 84 488
rect 43 411 83 413
rect 43 403 83 405
rect 135 379 175 381
rect -32 373 8 375
rect 135 371 175 373
rect -32 365 8 367
rect 40 339 80 341
rect 40 331 80 333
rect 40 253 80 255
rect 40 245 80 247
rect 132 221 172 223
rect -35 215 5 217
rect 132 213 172 215
rect -35 207 5 209
rect 37 181 77 183
rect 37 173 77 175
rect 37 49 77 51
rect 37 41 77 43
rect 129 17 169 19
rect -38 11 2 13
rect 129 9 169 11
rect -38 3 2 5
rect 34 -23 74 -21
rect 34 -31 74 -29
<< ptransistor >>
rect -12 722 28 724
rect -12 714 28 716
rect 80 690 120 692
rect -87 684 -47 686
rect 80 682 120 684
rect -87 676 -47 678
rect -15 650 25 652
rect -15 642 25 644
rect -15 566 25 568
rect -15 558 25 560
rect 77 534 117 536
rect -90 528 -50 530
rect 77 526 117 528
rect -90 520 -50 522
rect -18 494 22 496
rect -18 486 22 488
rect -19 411 21 413
rect -19 403 21 405
rect 73 379 113 381
rect -94 373 -54 375
rect 73 371 113 373
rect -94 365 -54 367
rect -22 339 18 341
rect -22 331 18 333
rect -22 253 18 255
rect -22 245 18 247
rect 70 221 110 223
rect -97 215 -57 217
rect 70 213 110 215
rect -97 207 -57 209
rect -25 181 15 183
rect -25 173 15 175
rect -25 49 15 51
rect -25 41 15 43
rect 67 17 107 19
rect -100 11 -60 13
rect 67 9 107 11
rect -100 3 -60 5
rect -28 -23 12 -21
rect -28 -31 12 -29
<< ndiffusion >>
rect 50 724 90 725
rect 50 721 90 722
rect 50 716 90 717
rect 50 713 90 714
rect 142 692 182 693
rect -25 686 15 687
rect -25 683 15 684
rect 142 689 182 690
rect 142 684 182 685
rect -25 678 15 679
rect 142 681 182 682
rect -25 675 15 676
rect 47 652 87 653
rect 47 649 87 650
rect 47 644 87 645
rect 47 641 87 642
rect 47 568 87 569
rect 47 565 87 566
rect 47 560 87 561
rect 47 557 87 558
rect 139 536 179 537
rect -28 530 12 531
rect -28 527 12 528
rect 139 533 179 534
rect 139 528 179 529
rect -28 522 12 523
rect 139 525 179 526
rect -28 519 12 520
rect 44 496 84 497
rect 44 493 84 494
rect 44 488 84 489
rect 44 485 84 486
rect 43 413 83 414
rect 43 410 83 411
rect 43 405 83 406
rect 43 402 83 403
rect 135 381 175 382
rect -32 375 8 376
rect -32 372 8 373
rect 135 378 175 379
rect 135 373 175 374
rect -32 367 8 368
rect 135 370 175 371
rect -32 364 8 365
rect 40 341 80 342
rect 40 338 80 339
rect 40 333 80 334
rect 40 330 80 331
rect 40 255 80 256
rect 40 252 80 253
rect 40 247 80 248
rect 40 244 80 245
rect 132 223 172 224
rect -35 217 5 218
rect -35 214 5 215
rect 132 220 172 221
rect 132 215 172 216
rect -35 209 5 210
rect 132 212 172 213
rect -35 206 5 207
rect 37 183 77 184
rect 37 180 77 181
rect 37 175 77 176
rect 37 172 77 173
rect 37 51 77 52
rect 37 48 77 49
rect 37 43 77 44
rect 37 40 77 41
rect 129 19 169 20
rect -38 13 2 14
rect -38 10 2 11
rect 129 16 169 17
rect 129 11 169 12
rect -38 5 2 6
rect 129 8 169 9
rect -38 2 2 3
rect 34 -21 74 -20
rect 34 -24 74 -23
rect 34 -29 74 -28
rect 34 -32 74 -31
<< pdiffusion >>
rect -12 724 28 725
rect -12 721 28 722
rect -12 716 28 717
rect -12 713 28 714
rect -87 686 -47 687
rect 80 692 120 693
rect 80 689 120 690
rect -87 683 -47 684
rect -87 678 -47 679
rect 80 684 120 685
rect 80 681 120 682
rect -87 675 -47 676
rect -15 652 25 653
rect -15 649 25 650
rect -15 644 25 645
rect -15 641 25 642
rect -15 568 25 569
rect -15 565 25 566
rect -15 560 25 561
rect -15 557 25 558
rect -90 530 -50 531
rect 77 536 117 537
rect 77 533 117 534
rect -90 527 -50 528
rect -90 522 -50 523
rect 77 528 117 529
rect 77 525 117 526
rect -90 519 -50 520
rect -18 496 22 497
rect -18 493 22 494
rect -18 488 22 489
rect -18 485 22 486
rect -19 413 21 414
rect -19 410 21 411
rect -19 405 21 406
rect -19 402 21 403
rect -94 375 -54 376
rect 73 381 113 382
rect 73 378 113 379
rect -94 372 -54 373
rect -94 367 -54 368
rect 73 373 113 374
rect 73 370 113 371
rect -94 364 -54 365
rect -22 341 18 342
rect -22 338 18 339
rect -22 333 18 334
rect -22 330 18 331
rect -22 255 18 256
rect -22 252 18 253
rect -22 247 18 248
rect -22 244 18 245
rect -97 217 -57 218
rect 70 223 110 224
rect 70 220 110 221
rect -97 214 -57 215
rect -97 209 -57 210
rect 70 215 110 216
rect 70 212 110 213
rect -97 206 -57 207
rect -25 183 15 184
rect -25 180 15 181
rect -25 175 15 176
rect -25 172 15 173
rect -25 51 15 52
rect -25 48 15 49
rect -25 43 15 44
rect -25 40 15 41
rect -100 13 -60 14
rect 67 19 107 20
rect 67 16 107 17
rect -100 10 -60 11
rect -100 5 -60 6
rect 67 11 107 12
rect 67 8 107 9
rect -100 2 -60 3
rect -28 -21 12 -20
rect -28 -24 12 -23
rect -28 -29 12 -28
rect -28 -32 12 -31
<< ndcontact >>
rect 50 725 90 729
rect 50 717 90 721
rect 50 709 90 713
rect -25 687 15 691
rect 142 693 182 697
rect -25 679 15 683
rect 142 685 182 689
rect 142 677 182 681
rect -25 671 15 675
rect 47 653 87 657
rect 47 645 87 649
rect 47 637 87 641
rect 47 569 87 573
rect 47 561 87 565
rect 47 553 87 557
rect -28 531 12 535
rect 139 537 179 541
rect -28 523 12 527
rect 139 529 179 533
rect 139 521 179 525
rect -28 515 12 519
rect 44 497 84 501
rect 44 489 84 493
rect 44 481 84 485
rect 43 414 83 418
rect 43 406 83 410
rect 43 398 83 402
rect -32 376 8 380
rect 135 382 175 386
rect -32 368 8 372
rect 135 374 175 378
rect 135 366 175 370
rect -32 360 8 364
rect 40 342 80 346
rect 40 334 80 338
rect 40 326 80 330
rect 40 256 80 260
rect 40 248 80 252
rect 40 240 80 244
rect -35 218 5 222
rect 132 224 172 228
rect -35 210 5 214
rect 132 216 172 220
rect 132 208 172 212
rect -35 202 5 206
rect 37 184 77 188
rect 37 176 77 180
rect 37 168 77 172
rect 37 52 77 56
rect 37 44 77 48
rect 37 36 77 40
rect -38 14 2 18
rect 129 20 169 24
rect -38 6 2 10
rect 129 12 169 16
rect 129 4 169 8
rect -38 -2 2 2
rect 34 -20 74 -16
rect 34 -28 74 -24
rect 34 -36 74 -32
<< pdcontact >>
rect -12 725 28 729
rect -12 717 28 721
rect -12 709 28 713
rect 80 693 120 697
rect -87 687 -47 691
rect 80 685 120 689
rect -87 679 -47 683
rect 80 677 120 681
rect -87 671 -47 675
rect -15 653 25 657
rect -15 645 25 649
rect -15 637 25 641
rect -15 569 25 573
rect -15 561 25 565
rect -15 553 25 557
rect 77 537 117 541
rect -90 531 -50 535
rect 77 529 117 533
rect -90 523 -50 527
rect 77 521 117 525
rect -90 515 -50 519
rect -18 497 22 501
rect -18 489 22 493
rect -18 481 22 485
rect -19 414 21 418
rect -19 406 21 410
rect -19 398 21 402
rect 73 382 113 386
rect -94 376 -54 380
rect 73 374 113 378
rect -94 368 -54 372
rect 73 366 113 370
rect -94 360 -54 364
rect -22 342 18 346
rect -22 334 18 338
rect -22 326 18 330
rect -22 256 18 260
rect -22 248 18 252
rect -22 240 18 244
rect 70 224 110 228
rect -97 218 -57 222
rect 70 216 110 220
rect -97 210 -57 214
rect 70 208 110 212
rect -97 202 -57 206
rect -25 184 15 188
rect -25 176 15 180
rect -25 168 15 172
rect -25 52 15 56
rect -25 44 15 48
rect -25 36 15 40
rect 67 20 107 24
rect -100 14 -60 18
rect 67 12 107 16
rect -100 6 -60 10
rect 67 4 107 8
rect -100 -2 -60 2
rect -28 -20 12 -16
rect -28 -28 12 -24
rect -28 -36 12 -32
<< polysilicon >>
rect -25 722 -12 724
rect 28 722 50 724
rect 90 722 93 724
rect -25 714 -12 716
rect 28 714 50 716
rect 90 714 93 716
rect 66 690 80 692
rect 120 690 142 692
rect 182 690 185 692
rect -100 684 -87 686
rect -47 684 -25 686
rect 15 684 18 686
rect 66 682 80 684
rect 120 682 142 684
rect 182 682 185 684
rect -100 676 -87 678
rect -47 676 -25 678
rect 15 676 18 678
rect -28 650 -15 652
rect 25 650 47 652
rect 87 650 90 652
rect -28 642 -15 644
rect 25 642 47 644
rect 87 642 90 644
rect -28 566 -15 568
rect 25 566 47 568
rect 87 566 90 568
rect -28 558 -15 560
rect 25 558 47 560
rect 87 558 90 560
rect 63 534 77 536
rect 117 534 139 536
rect 179 534 182 536
rect -103 528 -90 530
rect -50 528 -28 530
rect 12 528 15 530
rect 63 526 77 528
rect 117 526 139 528
rect 179 526 182 528
rect -103 520 -90 522
rect -50 520 -28 522
rect 12 520 15 522
rect -31 494 -18 496
rect 22 494 44 496
rect 84 494 87 496
rect -31 486 -18 488
rect 22 486 44 488
rect 84 486 87 488
rect -32 411 -19 413
rect 21 411 43 413
rect 83 411 86 413
rect -32 403 -19 405
rect 21 403 43 405
rect 83 403 86 405
rect 59 379 73 381
rect 113 379 135 381
rect 175 379 178 381
rect -107 373 -94 375
rect -54 373 -32 375
rect 8 373 11 375
rect 59 371 73 373
rect 113 371 135 373
rect 175 371 178 373
rect -107 365 -94 367
rect -54 365 -32 367
rect 8 365 11 367
rect -35 339 -22 341
rect 18 339 40 341
rect 80 339 83 341
rect -35 331 -22 333
rect 18 331 40 333
rect 80 331 83 333
rect -35 253 -22 255
rect 18 253 40 255
rect 80 253 83 255
rect -35 245 -22 247
rect 18 245 40 247
rect 80 245 83 247
rect 56 221 70 223
rect 110 221 132 223
rect 172 221 175 223
rect -110 215 -97 217
rect -57 215 -35 217
rect 5 215 8 217
rect 56 213 70 215
rect 110 213 132 215
rect 172 213 175 215
rect -110 207 -97 209
rect -57 207 -35 209
rect 5 207 8 209
rect -38 181 -25 183
rect 15 181 37 183
rect 77 181 80 183
rect -38 173 -25 175
rect 15 173 37 175
rect 77 173 80 175
rect -38 49 -25 51
rect 15 49 37 51
rect 77 49 80 51
rect -38 41 -25 43
rect 15 41 37 43
rect 77 41 80 43
rect 53 17 67 19
rect 107 17 129 19
rect 169 17 172 19
rect -113 11 -100 13
rect -60 11 -38 13
rect 2 11 5 13
rect 53 9 67 11
rect 107 9 129 11
rect 169 9 172 11
rect -113 3 -100 5
rect -60 3 -38 5
rect 2 3 5 5
rect -41 -23 -28 -21
rect 12 -23 34 -21
rect 74 -23 77 -21
rect -41 -31 -28 -29
rect 12 -31 34 -29
rect 74 -31 77 -29
<< polycontact >>
rect -29 721 -25 725
rect -29 713 -25 717
rect -104 683 -100 687
rect 62 689 66 693
rect -104 675 -100 679
rect 62 681 66 685
rect -32 649 -28 653
rect -32 641 -28 645
rect -32 565 -28 569
rect -32 557 -28 561
rect -107 527 -103 531
rect 59 533 63 537
rect -107 519 -103 523
rect 59 525 63 529
rect -35 493 -31 497
rect -35 485 -31 489
rect -36 410 -32 414
rect -36 402 -32 406
rect -111 372 -107 376
rect 55 378 59 382
rect -111 364 -107 368
rect 55 370 59 374
rect -39 338 -35 342
rect -39 330 -35 334
rect -39 252 -35 256
rect -39 244 -35 248
rect -114 214 -110 218
rect 52 220 56 224
rect -114 206 -110 210
rect 52 212 56 216
rect -42 180 -38 184
rect -42 172 -38 176
rect -42 48 -38 52
rect -42 40 -38 44
rect -117 10 -113 14
rect 49 16 53 20
rect -117 2 -113 6
rect 49 8 53 12
rect -45 -24 -41 -20
rect -45 -32 -41 -28
<< metal1 >>
rect -110 721 -29 725
rect -21 721 -17 750
rect 186 729 190 747
rect 28 725 36 729
rect 90 725 190 729
rect -110 689 -106 721
rect -21 717 -12 721
rect -35 713 -29 717
rect -110 688 -105 689
rect -127 687 -105 688
rect -47 687 -39 691
rect -127 683 -104 687
rect -110 682 -105 683
rect -96 679 -87 683
rect -110 677 -104 679
rect -125 675 -104 677
rect -125 672 -105 675
rect -109 645 -105 672
rect -96 668 -92 679
rect -43 675 -39 687
rect -34 675 -30 713
rect -21 702 -17 717
rect 32 713 36 725
rect 28 709 50 713
rect 39 693 43 709
rect 186 697 190 725
rect 15 687 23 691
rect 39 689 62 693
rect 70 689 74 697
rect 120 693 128 697
rect 182 693 190 697
rect 19 677 23 687
rect 70 685 80 689
rect 39 681 62 685
rect -47 671 -25 675
rect -38 670 -30 671
rect -38 653 -34 670
rect -38 649 -32 653
rect -24 649 -20 663
rect 25 653 33 657
rect -24 645 -15 649
rect -109 641 -32 645
rect -113 565 -32 569
rect -24 565 -20 645
rect 29 641 33 653
rect 39 641 43 681
rect 70 668 74 685
rect 124 681 128 693
rect 120 677 142 681
rect 132 670 136 677
rect 87 653 91 657
rect 186 657 190 693
rect 96 653 190 657
rect 25 637 47 641
rect 186 615 190 653
rect 183 610 190 615
rect 183 573 187 610
rect 25 569 33 573
rect 87 569 187 573
rect -113 533 -109 565
rect -24 561 -15 565
rect -38 557 -32 561
rect -113 532 -108 533
rect -130 531 -108 532
rect -50 531 -42 535
rect -130 527 -107 531
rect -113 526 -108 527
rect -99 523 -90 527
rect -113 521 -107 523
rect -128 519 -107 521
rect -128 516 -108 519
rect -112 489 -108 516
rect -99 512 -95 523
rect -46 519 -42 531
rect -37 519 -33 557
rect -24 546 -20 561
rect 29 557 33 569
rect 25 553 47 557
rect 36 537 40 553
rect 183 541 187 569
rect 12 531 20 535
rect 36 533 59 537
rect 67 533 71 541
rect 117 537 125 541
rect 179 537 187 541
rect 16 521 20 531
rect 67 529 77 533
rect 36 525 59 529
rect -50 515 -28 519
rect -41 514 -33 515
rect -41 497 -37 514
rect -41 493 -35 497
rect -27 493 -23 507
rect 22 497 30 501
rect -27 489 -18 493
rect -112 485 -35 489
rect -27 439 -23 489
rect 26 485 30 497
rect 36 485 40 525
rect 67 512 71 529
rect 121 525 125 537
rect 117 521 139 525
rect 129 514 133 521
rect 84 497 88 501
rect 183 501 187 537
rect 93 497 187 501
rect 22 481 44 485
rect 183 460 187 497
rect -28 434 -23 439
rect 179 454 187 460
rect 179 446 183 454
rect 179 434 184 446
rect -117 410 -36 414
rect -28 410 -24 434
rect 179 418 183 434
rect 21 414 29 418
rect 83 414 183 418
rect -117 378 -113 410
rect -28 406 -19 410
rect -42 402 -36 406
rect -117 377 -112 378
rect -134 376 -112 377
rect -54 376 -46 380
rect -134 372 -111 376
rect -117 371 -112 372
rect -103 368 -94 372
rect -117 366 -111 368
rect -132 364 -111 366
rect -132 361 -112 364
rect -116 334 -112 361
rect -103 357 -99 368
rect -50 364 -46 376
rect -41 364 -37 402
rect -28 391 -24 406
rect 25 402 29 414
rect 21 398 43 402
rect 32 382 36 398
rect 179 386 183 414
rect 8 376 16 380
rect 32 378 55 382
rect 63 378 67 386
rect 113 382 121 386
rect 175 382 183 386
rect 12 366 16 376
rect 63 374 73 378
rect 32 370 55 374
rect -54 360 -32 364
rect -45 359 -37 360
rect -45 342 -41 359
rect -45 338 -39 342
rect -31 338 -27 352
rect 18 342 26 346
rect -31 334 -22 338
rect -116 330 -39 334
rect -120 252 -39 256
rect -31 252 -27 334
rect 22 330 26 342
rect 32 330 36 370
rect 63 357 67 374
rect 117 370 121 382
rect 113 366 135 370
rect 125 359 129 366
rect 80 342 84 346
rect 179 346 183 382
rect 89 342 183 346
rect 18 326 40 330
rect 179 305 183 342
rect 176 299 183 305
rect 176 260 180 299
rect 18 256 26 260
rect 80 256 180 260
rect -120 220 -116 252
rect -31 248 -22 252
rect -45 244 -39 248
rect -120 219 -115 220
rect -137 218 -115 219
rect -57 218 -49 222
rect -137 214 -114 218
rect -120 213 -115 214
rect -106 210 -97 214
rect -120 208 -114 210
rect -135 206 -114 208
rect -135 203 -115 206
rect -119 176 -115 203
rect -106 199 -102 210
rect -53 206 -49 218
rect -44 206 -40 244
rect -31 233 -27 248
rect 22 244 26 256
rect 18 240 40 244
rect 29 224 33 240
rect 176 228 180 256
rect 5 218 13 222
rect 29 220 52 224
rect 60 220 64 228
rect 110 224 118 228
rect 172 224 180 228
rect 9 208 13 218
rect 60 216 70 220
rect 29 212 52 216
rect -57 202 -35 206
rect -48 201 -40 202
rect -48 184 -44 201
rect -48 180 -42 184
rect -34 180 -30 194
rect 15 184 23 188
rect -34 176 -25 180
rect -119 172 -42 176
rect -123 48 -42 52
rect -34 48 -30 176
rect 19 172 23 184
rect 29 172 33 212
rect 60 199 64 216
rect 114 212 118 224
rect 110 208 132 212
rect 122 201 126 208
rect 77 184 81 188
rect 176 188 180 224
rect 86 184 180 188
rect 15 168 37 172
rect 176 87 180 184
rect 172 83 180 87
rect 173 82 180 83
rect 173 56 177 82
rect 15 52 23 56
rect 77 52 177 56
rect -123 16 -119 48
rect -34 44 -25 48
rect -48 40 -42 44
rect -123 15 -118 16
rect -140 14 -118 15
rect -60 14 -52 18
rect -140 10 -117 14
rect -123 9 -118 10
rect -109 6 -100 10
rect -123 4 -117 6
rect -138 2 -117 4
rect -138 -1 -118 2
rect -122 -28 -118 -1
rect -109 -5 -105 6
rect -56 2 -52 14
rect -47 2 -43 40
rect -34 29 -30 44
rect 19 40 23 52
rect 15 36 37 40
rect 26 20 30 36
rect 173 24 177 52
rect 2 14 10 18
rect 26 16 49 20
rect 57 16 61 24
rect 107 20 115 24
rect 169 20 177 24
rect 6 4 10 14
rect 57 12 67 16
rect 26 8 49 12
rect -60 -2 -38 2
rect -51 -3 -43 -2
rect -51 -20 -47 -3
rect -51 -24 -45 -20
rect -37 -24 -33 -10
rect 12 -20 20 -16
rect -37 -28 -28 -24
rect -122 -32 -45 -28
rect -37 -80 -33 -28
rect 16 -32 20 -20
rect 26 -32 30 8
rect 57 -5 61 12
rect 111 8 115 20
rect 107 4 129 8
rect 119 -3 123 4
rect 74 -20 78 -16
rect 173 -16 177 20
rect 83 -20 177 -16
rect 12 -36 34 -32
rect 173 -63 177 -20
<< m2contact >>
rect -21 697 -16 702
rect 69 697 74 702
rect 19 672 24 677
rect -96 663 -91 668
rect -24 663 -19 668
rect 69 663 74 668
rect 132 665 137 670
rect 91 653 96 658
rect -24 541 -19 546
rect 66 541 71 546
rect 16 516 21 521
rect -99 507 -94 512
rect -27 507 -22 512
rect 66 507 71 512
rect 129 509 134 514
rect 88 497 93 502
rect -28 386 -23 391
rect 62 386 67 391
rect 12 361 17 366
rect -103 352 -98 357
rect -31 352 -26 357
rect 62 352 67 357
rect 125 354 130 359
rect 84 342 89 347
rect -31 228 -26 233
rect 59 228 64 233
rect 9 203 14 208
rect -106 194 -101 199
rect -34 194 -29 199
rect 59 194 64 199
rect 122 196 127 201
rect 81 184 86 189
rect -34 24 -29 29
rect 56 24 61 29
rect 6 -1 11 4
rect -109 -10 -104 -5
rect -37 -10 -32 -5
rect 56 -10 61 -5
rect 119 -8 124 -3
rect 78 -20 83 -15
<< metal2 >>
rect -16 697 69 702
rect 24 672 94 675
rect -91 663 -24 668
rect -19 663 69 668
rect 91 658 94 672
rect 132 646 136 665
rect 207 646 212 647
rect 132 642 212 646
rect -19 541 66 546
rect 21 516 91 519
rect -94 507 -27 512
rect -22 507 66 512
rect 88 502 91 516
rect 129 490 133 509
rect 204 490 209 491
rect 129 486 209 490
rect -23 386 62 391
rect 17 361 87 364
rect -98 352 -31 357
rect -26 352 62 357
rect 84 347 87 361
rect 125 335 129 354
rect 200 335 205 336
rect 125 331 205 335
rect -26 228 59 233
rect 14 203 84 206
rect -101 194 -34 199
rect -29 194 59 199
rect 81 189 84 203
rect 122 177 126 196
rect 197 177 202 178
rect 122 173 202 177
rect -29 24 56 29
rect 11 -1 81 2
rect -104 -10 -37 -5
rect -32 -10 56 -5
rect 78 -15 81 -1
rect 119 -27 123 -8
rect 194 -27 199 -26
rect 119 -31 199 -27
<< labels >>
rlabel metal1 -37 -80 -33 -76 1 vdd
rlabel metal1 173 -63 177 -59 1 gnd
rlabel metal2 194 -31 199 -26 1 p0
rlabel metal1 -140 10 -135 15 3 a0
rlabel metal1 -138 -1 -133 4 3 b0
rlabel metal1 -135 203 -130 208 1 b1
rlabel metal1 -137 214 -132 219 1 a1
rlabel metal1 -132 361 -127 366 1 b2
rlabel metal1 -134 372 -129 377 1 a2
rlabel metal1 -128 516 -123 521 1 b3
rlabel metal1 -130 527 -125 532 1 a3
rlabel metal1 -125 672 -120 677 1 b4
rlabel metal1 -127 683 -122 688 1 a4
rlabel metal2 207 642 212 647 7 p4
rlabel metal2 204 486 209 491 1 p3
rlabel metal2 200 331 205 336 1 p2
rlabel metal2 197 173 202 178 1 p1
<< end >>
