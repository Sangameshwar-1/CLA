magic
tech scmos
timestamp 1764137424
<< nwell >>
rect -226 1399 -174 1431
rect -225 1346 -169 1370
rect -216 1264 -164 1296
rect -216 1230 -160 1254
rect 483 1233 539 1257
rect -186 1140 -134 1172
rect -185 1110 -129 1134
rect 221 1032 273 1064
rect -737 971 -685 1003
rect -645 969 -593 971
rect 222 969 278 993
rect -812 933 -760 965
rect -646 937 -593 969
rect -740 899 -688 931
rect 39 865 91 944
rect -740 815 -688 847
rect -648 813 -596 815
rect -815 777 -763 809
rect -649 781 -596 813
rect 39 777 91 835
rect -743 743 -691 775
rect 39 715 91 765
rect 321 745 373 824
rect 894 722 946 754
rect 986 720 1038 722
rect -744 660 -692 692
rect 39 672 91 704
rect 819 684 871 716
rect 985 688 1038 720
rect -652 658 -600 660
rect -819 622 -767 654
rect -653 626 -600 658
rect 891 650 943 682
rect -747 588 -695 620
rect 891 566 943 598
rect 983 564 1035 566
rect -747 502 -695 534
rect -655 500 -603 502
rect 39 501 91 559
rect 816 528 868 560
rect 982 532 1035 564
rect -822 464 -770 496
rect -656 468 -603 500
rect -750 430 -698 462
rect 39 439 91 489
rect 276 438 328 496
rect 888 494 940 526
rect 39 396 91 428
rect 887 411 939 443
rect 979 409 1031 411
rect 812 373 864 405
rect 978 377 1031 409
rect 884 339 936 371
rect -750 298 -698 330
rect -658 296 -606 298
rect -825 260 -773 292
rect -659 264 -606 296
rect -753 226 -701 258
rect 39 223 91 273
rect 884 253 936 285
rect 976 251 1028 253
rect 39 173 91 205
rect 241 192 293 242
rect 809 215 861 247
rect 975 219 1028 251
rect 881 181 933 213
rect 40 30 92 62
rect 881 49 933 81
rect 973 47 1025 49
rect 214 11 266 43
rect 806 11 858 43
rect 972 15 1025 47
rect 878 -23 930 9
rect -679 -114 -627 -82
<< ntransistor >>
rect -158 1418 -118 1420
rect -158 1410 -118 1412
rect -161 1357 -141 1359
rect -148 1283 -108 1285
rect -148 1275 -108 1277
rect 547 1244 567 1246
rect -152 1241 -132 1243
rect -118 1159 -78 1161
rect -118 1151 -78 1153
rect -121 1121 -101 1123
rect 289 1051 329 1053
rect 289 1043 329 1045
rect -669 990 -629 992
rect -669 982 -629 984
rect 286 980 306 982
rect -577 958 -537 960
rect -744 952 -704 954
rect -577 950 -537 952
rect -744 944 -704 946
rect 107 928 207 930
rect -672 918 -632 920
rect -672 910 -632 912
rect 107 910 207 912
rect 107 902 207 904
rect 107 884 207 886
rect 107 876 207 878
rect -672 834 -632 836
rect -672 826 -632 828
rect 107 822 187 824
rect 107 814 187 816
rect 389 808 489 810
rect -580 802 -540 804
rect -747 796 -707 798
rect -580 794 -540 796
rect 107 796 187 798
rect -747 788 -707 790
rect 107 788 187 790
rect 389 790 489 792
rect 389 782 489 784
rect -675 762 -635 764
rect 389 764 489 766
rect -675 754 -635 756
rect 389 756 489 758
rect 107 752 167 754
rect 962 741 1002 743
rect 107 734 167 736
rect 962 733 1002 735
rect 107 726 167 728
rect 1054 709 1094 711
rect 887 703 927 705
rect 1054 701 1094 703
rect 887 695 927 697
rect 107 691 147 693
rect 107 683 147 685
rect -676 679 -636 681
rect -676 671 -636 673
rect 959 669 999 671
rect 959 661 999 663
rect -584 647 -544 649
rect -751 641 -711 643
rect -584 639 -544 641
rect -751 633 -711 635
rect -679 607 -639 609
rect -679 599 -639 601
rect 959 585 999 587
rect 959 577 999 579
rect 107 546 187 548
rect 1051 553 1091 555
rect 884 547 924 549
rect 107 538 187 540
rect 1051 545 1091 547
rect 884 539 924 541
rect -679 521 -639 523
rect 107 520 187 522
rect -679 513 -639 515
rect 107 512 187 514
rect 956 513 996 515
rect 956 505 996 507
rect -587 489 -547 491
rect -754 483 -714 485
rect -587 481 -547 483
rect -754 475 -714 477
rect 344 483 424 485
rect 107 476 167 478
rect 344 475 424 477
rect 107 458 167 460
rect -682 449 -642 451
rect 344 457 424 459
rect 107 450 167 452
rect 344 449 424 451
rect -682 441 -642 443
rect 955 430 995 432
rect 955 422 995 424
rect 107 415 147 417
rect 107 407 147 409
rect 1047 398 1087 400
rect 880 392 920 394
rect 1047 390 1087 392
rect 880 384 920 386
rect 952 358 992 360
rect 952 350 992 352
rect -682 317 -642 319
rect -682 309 -642 311
rect -590 285 -550 287
rect -757 279 -717 281
rect -590 277 -550 279
rect -757 271 -717 273
rect 952 272 992 274
rect 952 264 992 266
rect 107 260 167 262
rect -685 245 -645 247
rect 107 242 167 244
rect -685 237 -645 239
rect 107 234 167 236
rect 1044 240 1084 242
rect 877 234 917 236
rect 309 229 369 231
rect 1044 232 1084 234
rect 877 226 917 228
rect 309 211 369 213
rect 309 203 369 205
rect 949 200 989 202
rect 107 192 147 194
rect 949 192 989 194
rect 107 184 147 186
rect 949 68 989 70
rect 949 60 989 62
rect 108 49 148 51
rect 108 41 148 43
rect 282 30 322 32
rect 1041 36 1081 38
rect 874 30 914 32
rect 282 22 322 24
rect 1041 28 1081 30
rect 874 22 914 24
rect 946 -4 986 -2
rect 946 -12 986 -10
rect -611 -95 -571 -93
rect -611 -103 -571 -101
<< ptransistor >>
rect -220 1418 -180 1420
rect -220 1410 -180 1412
rect -215 1357 -175 1359
rect -210 1283 -170 1285
rect -210 1275 -170 1277
rect 493 1244 533 1246
rect -206 1241 -166 1243
rect -180 1159 -140 1161
rect -180 1151 -140 1153
rect -175 1121 -135 1123
rect 227 1051 267 1053
rect 227 1043 267 1045
rect -731 990 -691 992
rect -731 982 -691 984
rect 232 980 272 982
rect -639 958 -599 960
rect -806 952 -766 954
rect -639 950 -599 952
rect -806 944 -766 946
rect 45 928 85 930
rect -734 918 -694 920
rect -734 910 -694 912
rect 45 910 85 912
rect 45 902 85 904
rect 45 884 85 886
rect 45 876 85 878
rect -734 834 -694 836
rect -734 826 -694 828
rect 45 822 85 824
rect 45 814 85 816
rect 327 808 367 810
rect -642 802 -602 804
rect -809 796 -769 798
rect -642 794 -602 796
rect 45 796 85 798
rect -809 788 -769 790
rect 45 788 85 790
rect 327 790 367 792
rect 327 782 367 784
rect -737 762 -697 764
rect 327 764 367 766
rect -737 754 -697 756
rect 327 756 367 758
rect 45 752 85 754
rect 900 741 940 743
rect 45 734 85 736
rect 900 733 940 735
rect 45 726 85 728
rect 992 709 1032 711
rect 825 703 865 705
rect 992 701 1032 703
rect 825 695 865 697
rect 45 691 85 693
rect 45 683 85 685
rect -738 679 -698 681
rect -738 671 -698 673
rect 897 669 937 671
rect 897 661 937 663
rect -646 647 -606 649
rect -813 641 -773 643
rect -646 639 -606 641
rect -813 633 -773 635
rect -741 607 -701 609
rect -741 599 -701 601
rect 897 585 937 587
rect 897 577 937 579
rect 45 546 85 548
rect 989 553 1029 555
rect 822 547 862 549
rect 45 538 85 540
rect 989 545 1029 547
rect 822 539 862 541
rect -741 521 -701 523
rect 45 520 85 522
rect -741 513 -701 515
rect 45 512 85 514
rect 894 513 934 515
rect 894 505 934 507
rect -649 489 -609 491
rect -816 483 -776 485
rect -649 481 -609 483
rect -816 475 -776 477
rect 282 483 322 485
rect 45 476 85 478
rect 282 475 322 477
rect 45 458 85 460
rect -744 449 -704 451
rect 282 457 322 459
rect 45 450 85 452
rect 282 449 322 451
rect -744 441 -704 443
rect 893 430 933 432
rect 893 422 933 424
rect 45 415 85 417
rect 45 407 85 409
rect 985 398 1025 400
rect 818 392 858 394
rect 985 390 1025 392
rect 818 384 858 386
rect 890 358 930 360
rect 890 350 930 352
rect -744 317 -704 319
rect -744 309 -704 311
rect -652 285 -612 287
rect -819 279 -779 281
rect -652 277 -612 279
rect -819 271 -779 273
rect 890 272 930 274
rect 890 264 930 266
rect 45 260 85 262
rect -747 245 -707 247
rect 45 242 85 244
rect -747 237 -707 239
rect 45 234 85 236
rect 982 240 1022 242
rect 815 234 855 236
rect 247 229 287 231
rect 982 232 1022 234
rect 815 226 855 228
rect 247 211 287 213
rect 247 203 287 205
rect 887 200 927 202
rect 45 192 85 194
rect 887 192 927 194
rect 45 184 85 186
rect 887 68 927 70
rect 887 60 927 62
rect 46 49 86 51
rect 46 41 86 43
rect 220 30 260 32
rect 979 36 1019 38
rect 812 30 852 32
rect 220 22 260 24
rect 979 28 1019 30
rect 812 22 852 24
rect 884 -4 924 -2
rect 884 -12 924 -10
rect -673 -95 -633 -93
rect -673 -103 -633 -101
<< ndiffusion >>
rect -158 1420 -118 1421
rect -158 1417 -118 1418
rect -158 1412 -118 1413
rect -158 1409 -118 1410
rect -161 1359 -141 1360
rect -161 1356 -141 1357
rect -148 1285 -108 1286
rect -148 1282 -108 1283
rect -148 1277 -108 1278
rect -148 1274 -108 1275
rect 547 1246 567 1247
rect -152 1243 -132 1244
rect -152 1240 -132 1241
rect 547 1243 567 1244
rect -118 1161 -78 1162
rect -118 1158 -78 1159
rect -118 1153 -78 1154
rect -118 1150 -78 1151
rect -121 1123 -101 1124
rect -121 1120 -101 1121
rect 289 1053 329 1054
rect 289 1050 329 1051
rect 289 1045 329 1046
rect 289 1042 329 1043
rect -669 992 -629 993
rect -669 989 -629 990
rect -669 984 -629 985
rect 286 982 306 983
rect -669 981 -629 982
rect 286 979 306 980
rect -577 960 -537 961
rect -744 954 -704 955
rect -744 951 -704 952
rect -577 957 -537 958
rect -577 952 -537 953
rect -744 946 -704 947
rect -577 949 -537 950
rect -744 943 -704 944
rect 107 930 207 931
rect 107 927 207 928
rect -672 920 -632 921
rect -672 917 -632 918
rect -672 912 -632 913
rect -672 909 -632 910
rect 107 912 207 913
rect 107 909 207 910
rect 107 904 207 905
rect 107 901 207 902
rect 107 886 207 887
rect 107 883 207 884
rect 107 878 207 879
rect 107 875 207 876
rect -672 836 -632 837
rect -672 833 -632 834
rect -672 828 -632 829
rect -672 825 -632 826
rect 107 824 187 825
rect 107 821 187 822
rect 107 816 187 817
rect 107 813 187 814
rect 389 810 489 811
rect -580 804 -540 805
rect 389 807 489 808
rect -747 798 -707 799
rect -747 795 -707 796
rect -580 801 -540 802
rect -580 796 -540 797
rect 107 798 187 799
rect -747 790 -707 791
rect -580 793 -540 794
rect -747 787 -707 788
rect 107 795 187 796
rect 107 790 187 791
rect 389 792 489 793
rect 107 787 187 788
rect 389 789 489 790
rect 389 784 489 785
rect 389 781 489 782
rect -675 764 -635 765
rect 389 766 489 767
rect -675 761 -635 762
rect -675 756 -635 757
rect -675 753 -635 754
rect 389 763 489 764
rect 389 758 489 759
rect 107 754 167 755
rect 107 751 167 752
rect 389 755 489 756
rect 962 743 1002 744
rect 107 736 167 737
rect 107 733 167 734
rect 962 740 1002 741
rect 962 735 1002 736
rect 107 728 167 729
rect 962 732 1002 733
rect 107 725 167 726
rect 1054 711 1094 712
rect 887 705 927 706
rect 887 702 927 703
rect 1054 708 1094 709
rect 1054 703 1094 704
rect 887 697 927 698
rect 1054 700 1094 701
rect 107 693 147 694
rect 107 690 147 691
rect 887 694 927 695
rect 107 685 147 686
rect -676 681 -636 682
rect -676 678 -636 679
rect 107 682 147 683
rect -676 673 -636 674
rect -676 670 -636 671
rect 959 671 999 672
rect 959 668 999 669
rect 959 663 999 664
rect 959 660 999 661
rect -584 649 -544 650
rect -751 643 -711 644
rect -751 640 -711 641
rect -584 646 -544 647
rect -584 641 -544 642
rect -751 635 -711 636
rect -584 638 -544 639
rect -751 632 -711 633
rect -679 609 -639 610
rect -679 606 -639 607
rect -679 601 -639 602
rect -679 598 -639 599
rect 959 587 999 588
rect 959 584 999 585
rect 959 579 999 580
rect 959 576 999 577
rect 107 548 187 549
rect 1051 555 1091 556
rect 884 549 924 550
rect 107 545 187 546
rect 107 540 187 541
rect 884 546 924 547
rect 1051 552 1091 553
rect 1051 547 1091 548
rect 884 541 924 542
rect 1051 544 1091 545
rect 107 537 187 538
rect 884 538 924 539
rect -679 523 -639 524
rect -679 520 -639 521
rect 107 522 187 523
rect -679 515 -639 516
rect -679 512 -639 513
rect 107 519 187 520
rect 107 514 187 515
rect 956 515 996 516
rect 107 511 187 512
rect 956 512 996 513
rect 956 507 996 508
rect 956 504 996 505
rect -587 491 -547 492
rect -754 485 -714 486
rect -754 482 -714 483
rect -587 488 -547 489
rect -587 483 -547 484
rect -754 477 -714 478
rect -587 480 -547 481
rect 344 485 424 486
rect 107 478 167 479
rect -754 474 -714 475
rect 107 475 167 476
rect 344 482 424 483
rect 344 477 424 478
rect 344 474 424 475
rect 107 460 167 461
rect -682 451 -642 452
rect 107 457 167 458
rect 344 459 424 460
rect 107 452 167 453
rect -682 448 -642 449
rect 107 449 167 450
rect 344 456 424 457
rect 344 451 424 452
rect 344 448 424 449
rect -682 443 -642 444
rect -682 440 -642 441
rect 955 432 995 433
rect 955 429 995 430
rect 955 424 995 425
rect 107 417 147 418
rect 955 421 995 422
rect 107 414 147 415
rect 107 409 147 410
rect 107 406 147 407
rect 1047 400 1087 401
rect 880 394 920 395
rect 880 391 920 392
rect 1047 397 1087 398
rect 1047 392 1087 393
rect 880 386 920 387
rect 1047 389 1087 390
rect 880 383 920 384
rect 952 360 992 361
rect 952 357 992 358
rect 952 352 992 353
rect 952 349 992 350
rect -682 319 -642 320
rect -682 316 -642 317
rect -682 311 -642 312
rect -682 308 -642 309
rect -590 287 -550 288
rect -757 281 -717 282
rect -757 278 -717 279
rect -590 284 -550 285
rect -590 279 -550 280
rect -757 273 -717 274
rect -590 276 -550 277
rect 952 274 992 275
rect -757 270 -717 271
rect 952 271 992 272
rect 952 266 992 267
rect 107 262 167 263
rect 107 259 167 260
rect 952 263 992 264
rect -685 247 -645 248
rect -685 244 -645 245
rect 107 244 167 245
rect -685 239 -645 240
rect -685 236 -645 237
rect 107 241 167 242
rect 107 236 167 237
rect 107 233 167 234
rect 1044 242 1084 243
rect 877 236 917 237
rect 309 231 369 232
rect 309 228 369 229
rect 877 233 917 234
rect 1044 239 1084 240
rect 1044 234 1084 235
rect 877 228 917 229
rect 1044 231 1084 232
rect 877 225 917 226
rect 309 213 369 214
rect 309 210 369 211
rect 309 205 369 206
rect 309 202 369 203
rect 949 202 989 203
rect 107 194 147 195
rect 107 191 147 192
rect 949 199 989 200
rect 949 194 989 195
rect 949 191 989 192
rect 107 186 147 187
rect 107 183 147 184
rect 949 70 989 71
rect 949 67 989 68
rect 949 62 989 63
rect 949 59 989 60
rect 108 51 148 52
rect 108 48 148 49
rect 108 43 148 44
rect 108 40 148 41
rect 282 32 322 33
rect 282 29 322 30
rect 1041 38 1081 39
rect 874 32 914 33
rect 282 24 322 25
rect 282 21 322 22
rect 874 29 914 30
rect 1041 35 1081 36
rect 1041 30 1081 31
rect 874 24 914 25
rect 1041 27 1081 28
rect 874 21 914 22
rect 946 -2 986 -1
rect 946 -5 986 -4
rect 946 -10 986 -9
rect 946 -13 986 -12
rect -611 -93 -571 -92
rect -611 -96 -571 -95
rect -611 -101 -571 -100
rect -611 -104 -571 -103
<< pdiffusion >>
rect -220 1420 -180 1421
rect -220 1417 -180 1418
rect -220 1412 -180 1413
rect -220 1409 -180 1410
rect -215 1359 -175 1360
rect -215 1356 -175 1357
rect -210 1285 -170 1286
rect -210 1282 -170 1283
rect -210 1277 -170 1278
rect -210 1274 -170 1275
rect -206 1243 -166 1244
rect 493 1246 533 1247
rect 493 1243 533 1244
rect -206 1240 -166 1241
rect -180 1161 -140 1162
rect -180 1158 -140 1159
rect -180 1153 -140 1154
rect -180 1150 -140 1151
rect -175 1123 -135 1124
rect -175 1120 -135 1121
rect 227 1053 267 1054
rect 227 1050 267 1051
rect 227 1045 267 1046
rect 227 1042 267 1043
rect -731 992 -691 993
rect -731 989 -691 990
rect -731 984 -691 985
rect 232 982 272 983
rect -731 981 -691 982
rect 232 979 272 980
rect -806 954 -766 955
rect -639 960 -599 961
rect -639 957 -599 958
rect -806 951 -766 952
rect -806 946 -766 947
rect -639 952 -599 953
rect -639 949 -599 950
rect -806 943 -766 944
rect 45 930 85 931
rect 45 927 85 928
rect -734 920 -694 921
rect -734 917 -694 918
rect -734 912 -694 913
rect -734 909 -694 910
rect 45 912 85 913
rect 45 909 85 910
rect 45 904 85 905
rect 45 901 85 902
rect 45 886 85 887
rect 45 883 85 884
rect 45 878 85 879
rect 45 875 85 876
rect -734 836 -694 837
rect -734 833 -694 834
rect -734 828 -694 829
rect -734 825 -694 826
rect 45 824 85 825
rect 45 821 85 822
rect 45 816 85 817
rect 45 813 85 814
rect -809 798 -769 799
rect -642 804 -602 805
rect 327 810 367 811
rect 327 807 367 808
rect -642 801 -602 802
rect -809 795 -769 796
rect -809 790 -769 791
rect -642 796 -602 797
rect 45 798 85 799
rect 45 795 85 796
rect -642 793 -602 794
rect -809 787 -769 788
rect 45 790 85 791
rect 327 792 367 793
rect 327 789 367 790
rect 45 787 85 788
rect 327 784 367 785
rect 327 781 367 782
rect -737 764 -697 765
rect 327 766 367 767
rect 327 763 367 764
rect -737 761 -697 762
rect -737 756 -697 757
rect -737 753 -697 754
rect 45 754 85 755
rect 327 758 367 759
rect 327 755 367 756
rect 45 751 85 752
rect 45 736 85 737
rect 900 743 940 744
rect 900 740 940 741
rect 45 733 85 734
rect 45 728 85 729
rect 900 735 940 736
rect 900 732 940 733
rect 45 725 85 726
rect 825 705 865 706
rect 992 711 1032 712
rect 992 708 1032 709
rect 825 702 865 703
rect 45 693 85 694
rect 825 697 865 698
rect 992 703 1032 704
rect 992 700 1032 701
rect 825 694 865 695
rect 45 690 85 691
rect -738 681 -698 682
rect 45 685 85 686
rect 45 682 85 683
rect -738 678 -698 679
rect -738 673 -698 674
rect -738 670 -698 671
rect 897 671 937 672
rect 897 668 937 669
rect 897 663 937 664
rect 897 660 937 661
rect -813 643 -773 644
rect -646 649 -606 650
rect -646 646 -606 647
rect -813 640 -773 641
rect -813 635 -773 636
rect -646 641 -606 642
rect -646 638 -606 639
rect -813 632 -773 633
rect -741 609 -701 610
rect -741 606 -701 607
rect -741 601 -701 602
rect -741 598 -701 599
rect 897 587 937 588
rect 897 584 937 585
rect 897 579 937 580
rect 897 576 937 577
rect 45 548 85 549
rect 822 549 862 550
rect 989 555 1029 556
rect 989 552 1029 553
rect 822 546 862 547
rect 45 545 85 546
rect 45 540 85 541
rect 822 541 862 542
rect 989 547 1029 548
rect 989 544 1029 545
rect 822 538 862 539
rect 45 537 85 538
rect -741 523 -701 524
rect -741 520 -701 521
rect -741 515 -701 516
rect 45 522 85 523
rect 45 519 85 520
rect -741 512 -701 513
rect 45 514 85 515
rect 894 515 934 516
rect 894 512 934 513
rect 45 511 85 512
rect 894 507 934 508
rect 894 504 934 505
rect -816 485 -776 486
rect -649 491 -609 492
rect -649 488 -609 489
rect -816 482 -776 483
rect -816 477 -776 478
rect -649 483 -609 484
rect -649 480 -609 481
rect 45 478 85 479
rect 282 485 322 486
rect 282 482 322 483
rect 45 475 85 476
rect -816 474 -776 475
rect 282 477 322 478
rect 282 474 322 475
rect 45 460 85 461
rect 45 457 85 458
rect -744 451 -704 452
rect 45 452 85 453
rect 282 459 322 460
rect 282 456 322 457
rect 45 449 85 450
rect -744 448 -704 449
rect -744 443 -704 444
rect 282 451 322 452
rect 282 448 322 449
rect -744 440 -704 441
rect 893 432 933 433
rect 893 429 933 430
rect 45 417 85 418
rect 893 424 933 425
rect 893 421 933 422
rect 45 414 85 415
rect 45 409 85 410
rect 45 406 85 407
rect 818 394 858 395
rect 985 400 1025 401
rect 985 397 1025 398
rect 818 391 858 392
rect 818 386 858 387
rect 985 392 1025 393
rect 985 389 1025 390
rect 818 383 858 384
rect 890 360 930 361
rect 890 357 930 358
rect 890 352 930 353
rect 890 349 930 350
rect -744 319 -704 320
rect -744 316 -704 317
rect -744 311 -704 312
rect -744 308 -704 309
rect -819 281 -779 282
rect -652 287 -612 288
rect -652 284 -612 285
rect -819 278 -779 279
rect -819 273 -779 274
rect -652 279 -612 280
rect -652 276 -612 277
rect 890 274 930 275
rect 890 271 930 272
rect -819 270 -779 271
rect 45 262 85 263
rect 890 266 930 267
rect 890 263 930 264
rect 45 259 85 260
rect -747 247 -707 248
rect -747 244 -707 245
rect -747 239 -707 240
rect 45 244 85 245
rect 45 241 85 242
rect -747 236 -707 237
rect 45 236 85 237
rect 45 233 85 234
rect 247 231 287 232
rect 815 236 855 237
rect 982 242 1022 243
rect 982 239 1022 240
rect 815 233 855 234
rect 247 228 287 229
rect 815 228 855 229
rect 982 234 1022 235
rect 982 231 1022 232
rect 815 225 855 226
rect 247 213 287 214
rect 247 210 287 211
rect 247 205 287 206
rect 247 202 287 203
rect 45 194 85 195
rect 887 202 927 203
rect 887 199 927 200
rect 45 191 85 192
rect 45 186 85 187
rect 887 194 927 195
rect 887 191 927 192
rect 45 183 85 184
rect 887 70 927 71
rect 887 67 927 68
rect 887 62 927 63
rect 887 59 927 60
rect 46 51 86 52
rect 46 48 86 49
rect 46 43 86 44
rect 46 40 86 41
rect 220 32 260 33
rect 220 29 260 30
rect 220 24 260 25
rect 812 32 852 33
rect 979 38 1019 39
rect 979 35 1019 36
rect 812 29 852 30
rect 220 21 260 22
rect 812 24 852 25
rect 979 30 1019 31
rect 979 27 1019 28
rect 812 21 852 22
rect 884 -2 924 -1
rect 884 -5 924 -4
rect 884 -10 924 -9
rect 884 -13 924 -12
rect -673 -93 -633 -92
rect -673 -96 -633 -95
rect -673 -101 -633 -100
rect -673 -104 -633 -103
<< ndcontact >>
rect -158 1421 -118 1425
rect -158 1413 -118 1417
rect -158 1405 -118 1409
rect -161 1360 -141 1364
rect -161 1352 -141 1356
rect -148 1286 -108 1290
rect -148 1278 -108 1282
rect -148 1270 -108 1274
rect -152 1244 -132 1248
rect 547 1247 567 1251
rect -152 1236 -132 1240
rect 547 1239 567 1243
rect -118 1162 -78 1166
rect -118 1154 -78 1158
rect -118 1146 -78 1150
rect -121 1124 -101 1128
rect -121 1116 -101 1120
rect 289 1054 329 1058
rect 289 1046 329 1050
rect 289 1038 329 1042
rect -669 993 -629 997
rect -669 985 -629 989
rect 286 983 306 987
rect -669 977 -629 981
rect 286 975 306 979
rect -744 955 -704 959
rect -577 961 -537 965
rect -744 947 -704 951
rect -577 953 -537 957
rect -577 945 -537 949
rect -744 939 -704 943
rect 107 931 207 935
rect -672 921 -632 925
rect 107 923 207 927
rect -672 913 -632 917
rect 107 913 207 917
rect -672 905 -632 909
rect 107 905 207 909
rect 107 897 207 901
rect 107 887 207 891
rect 107 879 207 883
rect 107 871 207 875
rect -672 837 -632 841
rect -672 829 -632 833
rect -672 821 -632 825
rect 107 825 187 829
rect 107 817 187 821
rect 107 809 187 813
rect -747 799 -707 803
rect -580 805 -540 809
rect 389 811 489 815
rect 389 803 489 807
rect -747 791 -707 795
rect -580 797 -540 801
rect 107 799 187 803
rect -580 789 -540 793
rect 107 791 187 795
rect 389 793 489 797
rect -747 783 -707 787
rect 107 783 187 787
rect 389 785 489 789
rect 389 777 489 781
rect -675 765 -635 769
rect 389 767 489 771
rect -675 757 -635 761
rect -675 749 -635 753
rect 107 755 167 759
rect 389 759 489 763
rect 389 751 489 755
rect 107 747 167 751
rect 107 737 167 741
rect 962 744 1002 748
rect 107 729 167 733
rect 962 736 1002 740
rect 962 728 1002 732
rect 107 721 167 725
rect 887 706 927 710
rect 1054 712 1094 716
rect 107 694 147 698
rect 887 698 927 702
rect 1054 704 1094 708
rect 1054 696 1094 700
rect -676 682 -636 686
rect 887 690 927 694
rect 107 686 147 690
rect 107 678 147 682
rect -676 674 -636 678
rect -676 666 -636 670
rect 959 672 999 676
rect 959 664 999 668
rect 959 656 999 660
rect -751 644 -711 648
rect -584 650 -544 654
rect -751 636 -711 640
rect -584 642 -544 646
rect -584 634 -544 638
rect -751 628 -711 632
rect -679 610 -639 614
rect -679 602 -639 606
rect -679 594 -639 598
rect 959 588 999 592
rect 959 580 999 584
rect 959 572 999 576
rect 107 549 187 553
rect 884 550 924 554
rect 1051 556 1091 560
rect 107 541 187 545
rect 884 542 924 546
rect 1051 548 1091 552
rect 1051 540 1091 544
rect 107 533 187 537
rect 884 534 924 538
rect -679 524 -639 528
rect -679 516 -639 520
rect 107 523 187 527
rect -679 508 -639 512
rect 107 515 187 519
rect 956 516 996 520
rect 107 507 187 511
rect 956 508 996 512
rect 956 500 996 504
rect -754 486 -714 490
rect -587 492 -547 496
rect -754 478 -714 482
rect -587 484 -547 488
rect -587 476 -547 480
rect 107 479 167 483
rect 344 486 424 490
rect -754 470 -714 474
rect 107 471 167 475
rect 344 478 424 482
rect 344 470 424 474
rect 107 461 167 465
rect -682 452 -642 456
rect 107 453 167 457
rect 344 460 424 464
rect -682 444 -642 448
rect 107 445 167 449
rect 344 452 424 456
rect 344 444 424 448
rect -682 436 -642 440
rect 955 433 995 437
rect 107 418 147 422
rect 955 425 995 429
rect 955 417 995 421
rect 107 410 147 414
rect 107 402 147 406
rect 880 395 920 399
rect 1047 401 1087 405
rect 880 387 920 391
rect 1047 393 1087 397
rect 1047 385 1087 389
rect 880 379 920 383
rect 952 361 992 365
rect 952 353 992 357
rect 952 345 992 349
rect -682 320 -642 324
rect -682 312 -642 316
rect -682 304 -642 308
rect -757 282 -717 286
rect -590 288 -550 292
rect -757 274 -717 278
rect -590 280 -550 284
rect -590 272 -550 276
rect 952 275 992 279
rect -757 266 -717 270
rect 107 263 167 267
rect 952 267 992 271
rect 952 259 992 263
rect 107 255 167 259
rect -685 248 -645 252
rect -685 240 -645 244
rect 107 245 167 249
rect -685 232 -645 236
rect 107 237 167 241
rect 107 229 167 233
rect 309 232 369 236
rect 877 237 917 241
rect 1044 243 1084 247
rect 309 224 369 228
rect 877 229 917 233
rect 1044 235 1084 239
rect 1044 227 1084 231
rect 877 221 917 225
rect 309 214 369 218
rect 309 206 369 210
rect 107 195 147 199
rect 309 198 369 202
rect 949 203 989 207
rect 949 195 989 199
rect 107 187 147 191
rect 949 187 989 191
rect 107 179 147 183
rect 949 71 989 75
rect 949 63 989 67
rect 108 52 148 56
rect 949 55 989 59
rect 108 44 148 48
rect 108 36 148 40
rect 282 33 322 37
rect 874 33 914 37
rect 1041 39 1081 43
rect 282 25 322 29
rect 874 25 914 29
rect 1041 31 1081 35
rect 1041 23 1081 27
rect 282 17 322 21
rect 874 17 914 21
rect 946 -1 986 3
rect 946 -9 986 -5
rect 946 -17 986 -13
rect -611 -92 -571 -88
rect -611 -100 -571 -96
rect -611 -108 -571 -104
<< pdcontact >>
rect -220 1421 -180 1425
rect -220 1413 -180 1417
rect -220 1405 -180 1409
rect -215 1360 -175 1364
rect -215 1352 -175 1356
rect -210 1286 -170 1290
rect -210 1278 -170 1282
rect -210 1270 -170 1274
rect -206 1244 -166 1248
rect 493 1247 533 1251
rect -206 1236 -166 1240
rect 493 1239 533 1243
rect -180 1162 -140 1166
rect -180 1154 -140 1158
rect -180 1146 -140 1150
rect -175 1124 -135 1128
rect -175 1116 -135 1120
rect 227 1054 267 1058
rect 227 1046 267 1050
rect 227 1038 267 1042
rect -731 993 -691 997
rect -731 985 -691 989
rect 232 983 272 987
rect -731 977 -691 981
rect 232 975 272 979
rect -639 961 -599 965
rect -806 955 -766 959
rect -639 953 -599 957
rect -806 947 -766 951
rect -639 945 -599 949
rect -806 939 -766 943
rect 45 931 85 935
rect -734 921 -694 925
rect 45 923 85 927
rect -734 913 -694 917
rect 45 913 85 917
rect -734 905 -694 909
rect 45 905 85 909
rect 45 897 85 901
rect 45 887 85 891
rect 45 879 85 883
rect 45 871 85 875
rect -734 837 -694 841
rect -734 829 -694 833
rect -734 821 -694 825
rect 45 825 85 829
rect 45 817 85 821
rect 45 809 85 813
rect 327 811 367 815
rect -642 805 -602 809
rect -809 799 -769 803
rect 327 803 367 807
rect -642 797 -602 801
rect -809 791 -769 795
rect 45 799 85 803
rect -642 789 -602 793
rect 45 791 85 795
rect -809 783 -769 787
rect 327 793 367 797
rect 45 783 85 787
rect 327 785 367 789
rect 327 777 367 781
rect -737 765 -697 769
rect 327 767 367 771
rect -737 757 -697 761
rect 327 759 367 763
rect 45 755 85 759
rect -737 749 -697 753
rect 45 747 85 751
rect 327 751 367 755
rect 900 744 940 748
rect 45 737 85 741
rect 900 736 940 740
rect 45 729 85 733
rect 900 728 940 732
rect 45 721 85 725
rect 992 712 1032 716
rect 825 706 865 710
rect 992 704 1032 708
rect 825 698 865 702
rect 45 694 85 698
rect 992 696 1032 700
rect 45 686 85 690
rect -738 682 -698 686
rect 825 690 865 694
rect -738 674 -698 678
rect 45 678 85 682
rect 897 672 937 676
rect -738 666 -698 670
rect 897 664 937 668
rect 897 656 937 660
rect -646 650 -606 654
rect -813 644 -773 648
rect -646 642 -606 646
rect -813 636 -773 640
rect -646 634 -606 638
rect -813 628 -773 632
rect -741 610 -701 614
rect -741 602 -701 606
rect -741 594 -701 598
rect 897 588 937 592
rect 897 580 937 584
rect 897 572 937 576
rect 989 556 1029 560
rect 45 549 85 553
rect 822 550 862 554
rect 989 548 1029 552
rect 45 541 85 545
rect 822 542 862 546
rect 989 540 1029 544
rect 45 533 85 537
rect 822 534 862 538
rect -741 524 -701 528
rect 45 523 85 527
rect -741 516 -701 520
rect 45 515 85 519
rect -741 508 -701 512
rect 894 516 934 520
rect 45 507 85 511
rect 894 508 934 512
rect 894 500 934 504
rect -649 492 -609 496
rect -816 486 -776 490
rect -649 484 -609 488
rect -816 478 -776 482
rect 282 486 322 490
rect -649 476 -609 480
rect 45 479 85 483
rect 282 478 322 482
rect -816 470 -776 474
rect 45 471 85 475
rect 282 470 322 474
rect 45 461 85 465
rect 282 460 322 464
rect -744 452 -704 456
rect 45 453 85 457
rect 282 452 322 456
rect -744 444 -704 448
rect 45 445 85 449
rect 282 444 322 448
rect -744 436 -704 440
rect 893 433 933 437
rect 893 425 933 429
rect 45 418 85 422
rect 893 417 933 421
rect 45 410 85 414
rect 45 402 85 406
rect 985 401 1025 405
rect 818 395 858 399
rect 985 393 1025 397
rect 818 387 858 391
rect 985 385 1025 389
rect 818 379 858 383
rect 890 361 930 365
rect 890 353 930 357
rect 890 345 930 349
rect -744 320 -704 324
rect -744 312 -704 316
rect -744 304 -704 308
rect -652 288 -612 292
rect -819 282 -779 286
rect -652 280 -612 284
rect -819 274 -779 278
rect -652 272 -612 276
rect 890 275 930 279
rect -819 266 -779 270
rect 890 267 930 271
rect 45 263 85 267
rect 45 255 85 259
rect 890 259 930 263
rect -747 248 -707 252
rect 45 245 85 249
rect -747 240 -707 244
rect 982 243 1022 247
rect 45 237 85 241
rect -747 232 -707 236
rect 815 237 855 241
rect 45 229 85 233
rect 247 232 287 236
rect 982 235 1022 239
rect 815 229 855 233
rect 247 224 287 228
rect 982 227 1022 231
rect 815 221 855 225
rect 247 214 287 218
rect 247 206 287 210
rect 887 203 927 207
rect 45 195 85 199
rect 247 198 287 202
rect 887 195 927 199
rect 45 187 85 191
rect 887 187 927 191
rect 45 179 85 183
rect 887 71 927 75
rect 887 63 927 67
rect 46 52 86 56
rect 887 55 927 59
rect 46 44 86 48
rect 46 36 86 40
rect 979 39 1019 43
rect 220 33 260 37
rect 812 33 852 37
rect 220 25 260 29
rect 979 31 1019 35
rect 812 25 852 29
rect 220 17 260 21
rect 979 23 1019 27
rect 812 17 852 21
rect 884 -1 924 3
rect 884 -9 924 -5
rect 884 -17 924 -13
rect -673 -92 -633 -88
rect -673 -100 -633 -96
rect -673 -108 -633 -104
<< polysilicon >>
rect -233 1418 -220 1420
rect -180 1418 -158 1420
rect -118 1418 -115 1420
rect -233 1410 -220 1412
rect -180 1410 -158 1412
rect -118 1410 -115 1412
rect -168 1359 -164 1360
rect -218 1357 -215 1359
rect -175 1357 -161 1359
rect -141 1357 -138 1359
rect -223 1283 -210 1285
rect -170 1283 -148 1285
rect -108 1283 -105 1285
rect -223 1275 -210 1277
rect -170 1275 -148 1277
rect -108 1275 -105 1277
rect -159 1243 -155 1244
rect 540 1246 544 1247
rect 490 1244 493 1246
rect 533 1244 547 1246
rect 567 1244 570 1246
rect -209 1241 -206 1243
rect -166 1241 -152 1243
rect -132 1241 -129 1243
rect -193 1159 -180 1161
rect -140 1159 -118 1161
rect -78 1159 -75 1161
rect -193 1151 -180 1153
rect -140 1151 -118 1153
rect -78 1151 -75 1153
rect -128 1123 -124 1124
rect -178 1121 -175 1123
rect -135 1121 -121 1123
rect -101 1121 -98 1123
rect 214 1051 227 1053
rect 267 1051 289 1053
rect 329 1051 332 1053
rect 214 1043 227 1045
rect 267 1043 289 1045
rect 329 1043 332 1045
rect -744 990 -731 992
rect -691 990 -669 992
rect -629 990 -626 992
rect -744 982 -731 984
rect -691 982 -669 984
rect -629 982 -626 984
rect 279 982 283 983
rect 229 980 232 982
rect 272 980 286 982
rect 306 980 309 982
rect -653 958 -639 960
rect -599 958 -577 960
rect -537 958 -534 960
rect -819 952 -806 954
rect -766 952 -744 954
rect -704 952 -701 954
rect -653 950 -639 952
rect -599 950 -577 952
rect -537 950 -534 952
rect -819 944 -806 946
rect -766 944 -744 946
rect -704 944 -701 946
rect 32 928 45 930
rect 85 928 107 930
rect 207 928 210 930
rect -747 918 -734 920
rect -694 918 -672 920
rect -632 918 -629 920
rect -747 910 -734 912
rect -694 910 -672 912
rect -632 910 -629 912
rect 32 910 45 912
rect 85 910 107 912
rect 207 910 210 912
rect 32 902 45 904
rect 85 902 107 904
rect 207 902 210 904
rect 32 884 45 886
rect 85 884 107 886
rect 207 884 210 886
rect 32 876 45 878
rect 85 876 107 878
rect 207 876 210 878
rect -747 834 -734 836
rect -694 834 -672 836
rect -632 834 -629 836
rect -747 826 -734 828
rect -694 826 -672 828
rect -632 826 -629 828
rect 32 822 45 824
rect 85 822 107 824
rect 187 822 190 824
rect 32 814 45 816
rect 85 814 107 816
rect 187 814 190 816
rect 314 808 327 810
rect 367 808 389 810
rect 489 808 492 810
rect -656 802 -642 804
rect -602 802 -580 804
rect -540 802 -537 804
rect -822 796 -809 798
rect -769 796 -747 798
rect -707 796 -704 798
rect -656 794 -642 796
rect -602 794 -580 796
rect -540 794 -537 796
rect 32 796 45 798
rect 85 796 107 798
rect 187 796 190 798
rect -822 788 -809 790
rect -769 788 -747 790
rect -707 788 -704 790
rect 32 788 45 790
rect 85 788 107 790
rect 187 788 190 790
rect 314 790 327 792
rect 367 790 389 792
rect 489 790 492 792
rect 314 782 327 784
rect 367 782 389 784
rect 489 782 492 784
rect -750 762 -737 764
rect -697 762 -675 764
rect -635 762 -632 764
rect 314 764 327 766
rect 367 764 389 766
rect 489 764 492 766
rect -750 754 -737 756
rect -697 754 -675 756
rect -635 754 -632 756
rect 314 756 327 758
rect 367 756 389 758
rect 489 756 492 758
rect 32 752 45 754
rect 85 752 107 754
rect 167 752 170 754
rect 887 741 900 743
rect 940 741 962 743
rect 1002 741 1005 743
rect 32 734 45 736
rect 85 734 107 736
rect 167 734 170 736
rect 887 733 900 735
rect 940 733 962 735
rect 1002 733 1005 735
rect 32 726 45 728
rect 85 726 107 728
rect 167 726 170 728
rect 978 709 992 711
rect 1032 709 1054 711
rect 1094 709 1097 711
rect 812 703 825 705
rect 865 703 887 705
rect 927 703 930 705
rect 978 701 992 703
rect 1032 701 1054 703
rect 1094 701 1097 703
rect 812 695 825 697
rect 865 695 887 697
rect 927 695 930 697
rect 32 691 45 693
rect 85 691 107 693
rect 147 691 150 693
rect 32 683 45 685
rect 85 683 107 685
rect 147 683 150 685
rect -751 679 -738 681
rect -698 679 -676 681
rect -636 679 -633 681
rect -751 671 -738 673
rect -698 671 -676 673
rect -636 671 -633 673
rect 884 669 897 671
rect 937 669 959 671
rect 999 669 1002 671
rect 884 661 897 663
rect 937 661 959 663
rect 999 661 1002 663
rect -660 647 -646 649
rect -606 647 -584 649
rect -544 647 -541 649
rect -826 641 -813 643
rect -773 641 -751 643
rect -711 641 -708 643
rect -660 639 -646 641
rect -606 639 -584 641
rect -544 639 -541 641
rect -826 633 -813 635
rect -773 633 -751 635
rect -711 633 -708 635
rect -754 607 -741 609
rect -701 607 -679 609
rect -639 607 -636 609
rect -754 599 -741 601
rect -701 599 -679 601
rect -639 599 -636 601
rect 884 585 897 587
rect 937 585 959 587
rect 999 585 1002 587
rect 884 577 897 579
rect 937 577 959 579
rect 999 577 1002 579
rect 32 546 45 548
rect 85 546 107 548
rect 187 546 190 548
rect 975 553 989 555
rect 1029 553 1051 555
rect 1091 553 1094 555
rect 809 547 822 549
rect 862 547 884 549
rect 924 547 927 549
rect 32 538 45 540
rect 85 538 107 540
rect 187 538 190 540
rect 975 545 989 547
rect 1029 545 1051 547
rect 1091 545 1094 547
rect 809 539 822 541
rect 862 539 884 541
rect 924 539 927 541
rect -754 521 -741 523
rect -701 521 -679 523
rect -639 521 -636 523
rect 32 520 45 522
rect 85 520 107 522
rect 187 520 190 522
rect -754 513 -741 515
rect -701 513 -679 515
rect -639 513 -636 515
rect 32 512 45 514
rect 85 512 107 514
rect 187 512 190 514
rect 881 513 894 515
rect 934 513 956 515
rect 996 513 999 515
rect 881 505 894 507
rect 934 505 956 507
rect 996 505 999 507
rect -663 489 -649 491
rect -609 489 -587 491
rect -547 489 -544 491
rect -829 483 -816 485
rect -776 483 -754 485
rect -714 483 -711 485
rect -663 481 -649 483
rect -609 481 -587 483
rect -547 481 -544 483
rect -829 475 -816 477
rect -776 475 -754 477
rect -714 475 -711 477
rect 269 483 282 485
rect 322 483 344 485
rect 424 483 427 485
rect 32 476 45 478
rect 85 476 107 478
rect 167 476 170 478
rect 269 475 282 477
rect 322 475 344 477
rect 424 475 427 477
rect 32 458 45 460
rect 85 458 107 460
rect 167 458 170 460
rect -757 449 -744 451
rect -704 449 -682 451
rect -642 449 -639 451
rect 269 457 282 459
rect 322 457 344 459
rect 424 457 427 459
rect 32 450 45 452
rect 85 450 107 452
rect 167 450 170 452
rect 269 449 282 451
rect 322 449 344 451
rect 424 449 427 451
rect -757 441 -744 443
rect -704 441 -682 443
rect -642 441 -639 443
rect 880 430 893 432
rect 933 430 955 432
rect 995 430 998 432
rect 880 422 893 424
rect 933 422 955 424
rect 995 422 998 424
rect 32 415 45 417
rect 85 415 107 417
rect 147 415 150 417
rect 32 407 45 409
rect 85 407 107 409
rect 147 407 150 409
rect 971 398 985 400
rect 1025 398 1047 400
rect 1087 398 1090 400
rect 805 392 818 394
rect 858 392 880 394
rect 920 392 923 394
rect 971 390 985 392
rect 1025 390 1047 392
rect 1087 390 1090 392
rect 805 384 818 386
rect 858 384 880 386
rect 920 384 923 386
rect 877 358 890 360
rect 930 358 952 360
rect 992 358 995 360
rect 877 350 890 352
rect 930 350 952 352
rect 992 350 995 352
rect -757 317 -744 319
rect -704 317 -682 319
rect -642 317 -639 319
rect -757 309 -744 311
rect -704 309 -682 311
rect -642 309 -639 311
rect -666 285 -652 287
rect -612 285 -590 287
rect -550 285 -547 287
rect -832 279 -819 281
rect -779 279 -757 281
rect -717 279 -714 281
rect -666 277 -652 279
rect -612 277 -590 279
rect -550 277 -547 279
rect -832 271 -819 273
rect -779 271 -757 273
rect -717 271 -714 273
rect 877 272 890 274
rect 930 272 952 274
rect 992 272 995 274
rect 877 264 890 266
rect 930 264 952 266
rect 992 264 995 266
rect 32 260 45 262
rect 85 260 107 262
rect 167 260 170 262
rect -760 245 -747 247
rect -707 245 -685 247
rect -645 245 -642 247
rect 32 242 45 244
rect 85 242 107 244
rect 167 242 170 244
rect -760 237 -747 239
rect -707 237 -685 239
rect -645 237 -642 239
rect 32 234 45 236
rect 85 234 107 236
rect 167 234 170 236
rect 968 240 982 242
rect 1022 240 1044 242
rect 1084 240 1087 242
rect 802 234 815 236
rect 855 234 877 236
rect 917 234 920 236
rect 234 229 247 231
rect 287 229 309 231
rect 369 229 372 231
rect 968 232 982 234
rect 1022 232 1044 234
rect 1084 232 1087 234
rect 802 226 815 228
rect 855 226 877 228
rect 917 226 920 228
rect 234 211 247 213
rect 287 211 309 213
rect 369 211 372 213
rect 234 203 247 205
rect 287 203 309 205
rect 369 203 372 205
rect 874 200 887 202
rect 927 200 949 202
rect 989 200 992 202
rect 32 192 45 194
rect 85 192 107 194
rect 147 192 150 194
rect 874 192 887 194
rect 927 192 949 194
rect 989 192 992 194
rect 32 184 45 186
rect 85 184 107 186
rect 147 184 150 186
rect 874 68 887 70
rect 927 68 949 70
rect 989 68 992 70
rect 874 60 887 62
rect 927 60 949 62
rect 989 60 992 62
rect 33 49 46 51
rect 86 49 108 51
rect 148 49 151 51
rect 33 41 46 43
rect 86 41 108 43
rect 148 41 151 43
rect 207 30 220 32
rect 260 30 282 32
rect 322 30 325 32
rect 965 36 979 38
rect 1019 36 1041 38
rect 1081 36 1084 38
rect 799 30 812 32
rect 852 30 874 32
rect 914 30 917 32
rect 207 22 220 24
rect 260 22 282 24
rect 322 22 325 24
rect 965 28 979 30
rect 1019 28 1041 30
rect 1081 28 1084 30
rect 799 22 812 24
rect 852 22 874 24
rect 914 22 917 24
rect 871 -4 884 -2
rect 924 -4 946 -2
rect 986 -4 989 -2
rect 871 -12 884 -10
rect 924 -12 946 -10
rect 986 -12 989 -10
rect -686 -95 -673 -93
rect -633 -95 -611 -93
rect -571 -95 -568 -93
rect -686 -103 -673 -101
rect -633 -103 -611 -101
rect -571 -103 -568 -101
<< polycontact >>
rect -237 1417 -233 1421
rect -237 1409 -233 1413
rect -168 1360 -164 1364
rect -227 1282 -223 1286
rect -227 1274 -223 1278
rect -159 1244 -155 1248
rect 540 1247 544 1251
rect -197 1158 -193 1162
rect -197 1150 -193 1154
rect -128 1124 -124 1128
rect 210 1050 214 1054
rect 210 1042 214 1046
rect -748 989 -744 993
rect -748 981 -744 985
rect 279 983 283 987
rect -823 951 -819 955
rect -657 957 -653 961
rect -823 943 -819 947
rect -657 949 -653 953
rect 28 927 32 931
rect -751 917 -747 921
rect -751 909 -747 913
rect 28 909 32 913
rect 28 901 32 905
rect 28 883 32 887
rect 28 875 32 879
rect -751 833 -747 837
rect -751 825 -747 829
rect 28 821 32 825
rect 28 813 32 817
rect -826 795 -822 799
rect -660 801 -656 805
rect 310 807 314 811
rect -826 787 -822 791
rect -660 793 -656 797
rect 28 795 32 799
rect 28 787 32 791
rect 310 789 314 793
rect 310 781 314 785
rect -754 761 -750 765
rect 310 763 314 767
rect -754 753 -750 757
rect 28 751 32 755
rect 310 755 314 759
rect 28 733 32 737
rect 883 740 887 744
rect 28 725 32 729
rect 883 732 887 736
rect 808 702 812 706
rect 974 708 978 712
rect 28 690 32 694
rect 808 694 812 698
rect 974 700 978 704
rect -755 678 -751 682
rect 28 682 32 686
rect -755 670 -751 674
rect 880 668 884 672
rect 880 660 884 664
rect -830 640 -826 644
rect -664 646 -660 650
rect -830 632 -826 636
rect -664 638 -660 642
rect -758 606 -754 610
rect -758 598 -754 602
rect 880 584 884 588
rect 880 576 884 580
rect 28 545 32 549
rect 805 546 809 550
rect 971 552 975 556
rect 28 537 32 541
rect 805 538 809 542
rect 971 544 975 548
rect -758 520 -754 524
rect -758 512 -754 516
rect 28 519 32 523
rect 28 511 32 515
rect 877 512 881 516
rect 877 504 881 508
rect -833 482 -829 486
rect -667 488 -663 492
rect -833 474 -829 478
rect -667 480 -663 484
rect 28 475 32 479
rect 265 482 269 486
rect 265 474 269 478
rect 28 457 32 461
rect -761 448 -757 452
rect 28 449 32 453
rect 265 456 269 460
rect -761 440 -757 444
rect 265 448 269 452
rect 876 429 880 433
rect 28 414 32 418
rect 876 421 880 425
rect 28 406 32 410
rect 801 391 805 395
rect 967 397 971 401
rect 801 383 805 387
rect 967 389 971 393
rect 873 357 877 361
rect 873 349 877 353
rect -761 316 -757 320
rect -761 308 -757 312
rect -836 278 -832 282
rect -670 284 -666 288
rect -836 270 -832 274
rect -670 276 -666 280
rect 873 271 877 275
rect 28 259 32 263
rect 873 263 877 267
rect -764 244 -760 248
rect -764 236 -760 240
rect 28 241 32 245
rect 28 233 32 237
rect 230 228 234 232
rect 798 233 802 237
rect 964 239 968 243
rect 798 225 802 229
rect 964 231 968 235
rect 230 210 234 214
rect 230 202 234 206
rect 28 191 32 195
rect 870 199 874 203
rect 28 183 32 187
rect 870 191 874 195
rect 870 67 874 71
rect 870 59 874 63
rect 29 48 33 52
rect 29 40 33 44
rect 203 29 207 33
rect 203 21 207 25
rect 795 29 799 33
rect 961 35 965 39
rect 795 21 799 25
rect 961 27 965 31
rect 867 -5 871 -1
rect 867 -13 871 -9
rect -690 -96 -686 -92
rect -690 -104 -686 -100
<< metal1 >>
rect -180 1421 -172 1425
rect -118 1421 -110 1425
rect -947 1417 -237 1421
rect -947 476 -943 1417
rect -229 1413 -220 1417
rect -934 1409 -237 1413
rect -176 1409 -172 1421
rect -934 1021 -930 1409
rect -180 1405 -158 1409
rect -168 1403 -163 1405
rect -225 1364 -221 1370
rect -168 1364 -164 1403
rect -137 1364 -133 1370
rect -225 1360 -215 1364
rect -141 1360 -133 1364
rect -225 1346 -221 1360
rect -168 1356 -164 1360
rect -175 1352 -161 1356
rect -168 1310 -164 1352
rect -137 1346 -133 1360
rect -170 1286 -162 1290
rect -108 1286 -100 1290
rect -936 1011 -930 1021
rect -924 1282 -227 1286
rect -936 487 -931 1011
rect -924 668 -920 1282
rect -219 1278 -210 1282
rect -913 1274 -227 1278
rect -166 1274 -162 1286
rect -913 699 -909 1274
rect -170 1270 -148 1274
rect -216 1248 -212 1254
rect -159 1248 -155 1270
rect -128 1248 -124 1254
rect -216 1244 -206 1248
rect -132 1244 -124 1248
rect -216 1230 -212 1244
rect -166 1236 -152 1240
rect -159 1221 -155 1236
rect -128 1230 -124 1244
rect 483 1251 487 1257
rect 540 1251 544 1267
rect 571 1251 575 1257
rect 483 1247 493 1251
rect 567 1247 575 1251
rect 483 1233 487 1247
rect 540 1243 544 1247
rect 533 1239 547 1243
rect 540 1229 544 1239
rect 571 1233 575 1247
rect -140 1162 -132 1166
rect -78 1162 -70 1166
rect -901 1158 -197 1162
rect -901 788 -897 1158
rect -189 1154 -180 1158
rect -887 1150 -197 1154
rect -136 1150 -132 1162
rect -887 800 -883 1150
rect -140 1146 -118 1150
rect -185 1128 -181 1134
rect -128 1128 -124 1146
rect -97 1128 -93 1134
rect -185 1124 -175 1128
rect -101 1124 -93 1128
rect -185 1110 -181 1124
rect -135 1116 -121 1120
rect -128 1112 -124 1116
rect -97 1110 -93 1124
rect -872 1054 208 1058
rect 267 1054 275 1058
rect 329 1054 337 1058
rect -872 1053 210 1054
rect -872 945 -867 1053
rect 204 1050 210 1053
rect 218 1046 227 1050
rect -860 1042 210 1046
rect 271 1042 275 1054
rect -860 1039 -856 1042
rect -860 1029 -854 1039
rect 267 1038 289 1042
rect -859 956 -854 1029
rect -829 989 -748 993
rect -740 989 -736 1018
rect -533 997 -529 1015
rect -691 993 -683 997
rect -629 993 -529 997
rect 279 1011 283 1038
rect 279 1007 295 1011
rect -829 957 -825 989
rect -740 985 -731 989
rect -754 981 -748 985
rect -829 956 -824 957
rect -859 955 -824 956
rect -766 955 -758 959
rect -859 951 -823 955
rect -829 950 -824 951
rect -815 947 -806 951
rect -829 945 -823 947
rect -872 943 -823 945
rect -872 940 -824 943
rect -828 913 -824 940
rect -815 936 -811 947
rect -762 943 -758 955
rect -753 943 -749 981
rect -740 970 -736 985
rect -687 981 -683 993
rect -691 977 -669 981
rect -680 961 -676 977
rect -533 965 -529 993
rect 222 987 226 993
rect 279 987 283 1007
rect 310 987 314 993
rect 222 983 232 987
rect 306 983 314 987
rect 222 969 226 983
rect 279 979 283 983
rect 272 975 286 979
rect -704 955 -696 959
rect -680 957 -657 961
rect -649 957 -645 965
rect -599 961 -591 965
rect -537 961 -529 965
rect -700 945 -696 955
rect -649 953 -639 957
rect -680 949 -657 953
rect -766 939 -744 943
rect -757 938 -749 939
rect -757 921 -753 938
rect -757 917 -751 921
rect -743 917 -739 931
rect -694 921 -686 925
rect -743 913 -734 917
rect -828 909 -751 913
rect -832 833 -751 837
rect -743 833 -739 913
rect -690 909 -686 921
rect -680 909 -676 949
rect -649 936 -645 953
rect -595 949 -591 961
rect -599 945 -577 949
rect -587 938 -583 945
rect -632 921 -628 925
rect -533 925 -529 961
rect -1 927 0 931
rect 5 927 28 931
rect 37 927 41 952
rect 85 931 93 935
rect 207 931 215 935
rect -623 921 -529 925
rect 36 923 45 927
rect -694 905 -672 909
rect -533 883 -529 921
rect -536 878 -529 883
rect -231 887 -227 914
rect 11 909 28 913
rect 37 909 41 923
rect 89 917 93 931
rect 279 929 283 975
rect 310 969 314 983
rect 85 913 93 917
rect 101 923 107 927
rect 101 917 105 923
rect 101 913 107 917
rect 36 905 45 909
rect -209 901 28 905
rect -231 883 28 887
rect 37 883 41 905
rect 89 901 93 913
rect 85 897 94 901
rect 101 897 107 901
rect 89 891 93 897
rect 85 887 93 891
rect 101 891 105 897
rect 101 887 107 891
rect -536 841 -532 878
rect -694 837 -686 841
rect -632 837 -532 841
rect -832 801 -828 833
rect -743 829 -734 833
rect -757 825 -751 829
rect -832 800 -827 801
rect -887 799 -827 800
rect -769 799 -761 803
rect -887 796 -826 799
rect -849 795 -826 796
rect -832 794 -827 795
rect -818 791 -809 795
rect -832 789 -826 791
rect -847 788 -826 789
rect -901 787 -826 788
rect -901 784 -827 787
rect -831 757 -827 784
rect -818 780 -814 791
rect -765 787 -761 799
rect -756 787 -752 825
rect -743 814 -739 829
rect -690 825 -686 837
rect -694 821 -672 825
rect -683 805 -679 821
rect -536 809 -532 837
rect -707 799 -699 803
rect -683 801 -660 805
rect -652 801 -648 809
rect -602 805 -594 809
rect -540 805 -532 809
rect -703 789 -699 799
rect -652 797 -642 801
rect -683 793 -660 797
rect -769 783 -747 787
rect -760 782 -752 783
rect -760 765 -756 782
rect -760 761 -754 765
rect -746 761 -742 775
rect -697 765 -689 769
rect -746 757 -737 761
rect -831 753 -754 757
rect -746 707 -742 757
rect -693 753 -689 765
rect -683 753 -679 793
rect -652 780 -648 797
rect -598 793 -594 805
rect -602 789 -580 793
rect -590 782 -586 789
rect -635 765 -631 769
rect -536 769 -532 805
rect -626 765 -532 769
rect -697 749 -675 753
rect -536 728 -532 765
rect -747 702 -742 707
rect -540 722 -532 728
rect -540 714 -536 722
rect -540 702 -535 714
rect -924 663 -918 668
rect -913 667 -906 699
rect -923 634 -918 663
rect -911 645 -906 667
rect -836 678 -755 682
rect -747 678 -743 702
rect -540 686 -536 702
rect -698 682 -690 686
rect -636 682 -536 686
rect -836 646 -832 678
rect -747 674 -738 678
rect -761 670 -755 674
rect -836 645 -831 646
rect -911 644 -831 645
rect -773 644 -765 648
rect -911 640 -830 644
rect -836 639 -831 640
rect -822 636 -813 640
rect -836 634 -830 636
rect -923 632 -830 634
rect -923 629 -831 632
rect -835 602 -831 629
rect -822 625 -818 636
rect -769 632 -765 644
rect -760 632 -756 670
rect -747 659 -743 674
rect -694 670 -690 682
rect -698 666 -676 670
rect -687 650 -683 666
rect -540 654 -536 682
rect -711 644 -703 648
rect -687 646 -664 650
rect -656 646 -652 654
rect -606 650 -598 654
rect -544 650 -536 654
rect -707 634 -703 644
rect -656 642 -646 646
rect -687 638 -664 642
rect -773 628 -751 632
rect -764 627 -756 628
rect -764 610 -760 627
rect -764 606 -758 610
rect -750 606 -746 620
rect -701 610 -693 614
rect -750 602 -741 606
rect -835 598 -758 602
rect -839 520 -758 524
rect -750 520 -746 602
rect -697 598 -693 610
rect -687 598 -683 638
rect -656 625 -652 642
rect -602 638 -598 650
rect -606 634 -584 638
rect -594 627 -590 634
rect -639 610 -635 614
rect -540 614 -536 650
rect -630 610 -536 614
rect -701 594 -679 598
rect -540 573 -536 610
rect -543 567 -536 573
rect -543 528 -539 567
rect -701 524 -693 528
rect -639 524 -539 528
rect -839 488 -835 520
rect -750 516 -741 520
rect -764 512 -758 516
rect -839 487 -834 488
rect -936 486 -834 487
rect -776 486 -768 490
rect -936 482 -833 486
rect -839 481 -834 482
rect -825 478 -816 482
rect -839 476 -833 478
rect -947 474 -833 476
rect -946 471 -834 474
rect -838 444 -834 471
rect -825 467 -821 478
rect -772 474 -768 486
rect -763 474 -759 512
rect -750 501 -746 516
rect -697 512 -693 524
rect -701 508 -679 512
rect -690 492 -686 508
rect -543 496 -539 524
rect -714 486 -706 490
rect -690 488 -667 492
rect -659 488 -655 496
rect -609 492 -601 496
rect -547 492 -539 496
rect -710 476 -706 486
rect -659 484 -649 488
rect -690 480 -667 484
rect -776 470 -754 474
rect -767 469 -759 470
rect -767 452 -763 469
rect -767 448 -761 452
rect -753 448 -749 462
rect -704 452 -696 456
rect -753 444 -744 448
rect -838 440 -761 444
rect -842 316 -761 320
rect -753 316 -749 444
rect -700 440 -696 452
rect -690 440 -686 480
rect -659 467 -655 484
rect -605 480 -601 492
rect -609 476 -587 480
rect -597 469 -593 476
rect -642 452 -638 456
rect -543 456 -539 492
rect -633 452 -539 456
rect -704 436 -682 440
rect -543 355 -539 452
rect -547 351 -539 355
rect -546 350 -539 351
rect -231 523 -227 883
rect 36 879 45 883
rect 15 875 28 879
rect -2 821 28 825
rect 37 821 41 879
rect 89 875 93 887
rect 85 871 107 875
rect 97 859 101 871
rect 97 855 304 859
rect 85 825 93 829
rect 187 825 195 829
rect 36 817 45 821
rect 8 813 28 817
rect -214 795 28 799
rect 37 795 41 817
rect 89 813 93 825
rect 85 809 94 813
rect 101 809 107 813
rect 300 811 304 855
rect 89 803 93 809
rect 85 799 93 803
rect 101 803 105 809
rect 300 807 310 811
rect 317 807 321 824
rect 367 811 375 815
rect 489 811 497 815
rect 300 806 304 807
rect 317 803 327 807
rect 101 799 107 803
rect 36 791 45 795
rect 15 787 28 791
rect 37 759 41 791
rect 89 787 93 799
rect 212 789 310 793
rect 317 789 321 803
rect 371 797 375 811
rect 367 793 375 797
rect 383 803 389 807
rect 383 797 387 803
rect 383 793 389 797
rect 85 783 107 787
rect 97 778 101 783
rect 212 778 216 789
rect 317 785 327 789
rect 97 774 216 778
rect 231 781 310 785
rect 36 755 45 759
rect 167 755 174 759
rect 3 751 28 755
rect 6 733 28 737
rect 37 733 41 755
rect 85 747 93 751
rect 89 741 93 747
rect 85 737 93 741
rect 101 747 107 751
rect 101 741 105 747
rect 101 737 107 741
rect 36 729 45 733
rect 15 725 28 729
rect 11 690 28 694
rect 37 690 41 729
rect 89 725 93 737
rect 85 721 107 725
rect 100 716 104 721
rect 231 716 235 781
rect 100 712 235 716
rect 244 763 310 767
rect 317 763 321 785
rect 371 781 375 793
rect 367 777 376 781
rect 383 777 389 781
rect 371 771 375 777
rect 367 767 375 771
rect 383 771 387 777
rect 383 767 389 771
rect 85 694 93 698
rect 147 694 155 698
rect 36 686 45 690
rect -18 682 28 686
rect -18 646 -14 682
rect 37 658 41 686
rect 89 682 93 694
rect 85 678 107 682
rect 100 673 104 678
rect 244 673 248 763
rect 317 759 327 763
rect 300 755 310 759
rect 100 669 248 673
rect 317 658 321 759
rect 371 755 375 767
rect 367 751 389 755
rect 379 709 383 751
rect 802 740 883 744
rect 891 740 895 769
rect 1098 748 1102 766
rect 940 744 948 748
rect 1002 744 1102 748
rect 379 707 575 709
rect 802 708 806 740
rect 891 736 900 740
rect 877 732 883 736
rect 802 707 807 708
rect 379 706 807 707
rect 865 706 873 710
rect 379 705 808 706
rect 571 702 808 705
rect 571 698 575 702
rect 802 701 807 702
rect 816 698 825 702
rect 802 696 808 698
rect 787 694 808 696
rect 787 691 807 694
rect 803 664 807 691
rect 816 687 820 698
rect 869 694 873 706
rect 878 694 882 732
rect 891 721 895 736
rect 944 732 948 744
rect 940 728 962 732
rect 951 712 955 728
rect 1098 716 1102 744
rect 927 706 935 710
rect 951 708 974 712
rect 982 708 986 716
rect 1032 712 1040 716
rect 1094 712 1102 716
rect 931 696 935 706
rect 982 704 992 708
rect 951 700 974 704
rect 865 690 887 694
rect 874 689 882 690
rect 874 672 878 689
rect 874 668 880 672
rect 888 668 892 682
rect 937 672 945 676
rect 888 664 897 668
rect 803 660 880 664
rect 37 654 321 658
rect 37 646 41 654
rect -18 642 269 646
rect -8 545 28 549
rect 37 545 41 642
rect 799 584 880 588
rect 888 584 892 664
rect 941 660 945 672
rect 951 660 955 700
rect 982 687 986 704
rect 1036 700 1040 712
rect 1032 696 1054 700
rect 1044 689 1048 696
rect 999 672 1003 676
rect 1098 676 1102 712
rect 1008 672 1102 676
rect 937 656 959 660
rect 1098 634 1102 672
rect 1095 629 1102 634
rect 1095 592 1099 629
rect 937 588 945 592
rect 999 588 1099 592
rect 85 549 93 553
rect 187 549 195 553
rect 799 552 803 584
rect 888 580 897 584
rect 874 576 880 580
rect 799 551 804 552
rect 546 550 804 551
rect 862 550 870 554
rect 36 541 45 545
rect -209 537 28 541
rect -231 519 28 523
rect 37 519 41 541
rect 89 537 93 549
rect 546 546 805 550
rect 85 533 94 537
rect 101 533 107 537
rect 89 527 93 533
rect 85 523 93 527
rect 101 527 105 533
rect 101 523 107 527
rect -231 446 -227 519
rect 36 515 45 519
rect 12 511 28 515
rect 37 483 41 515
rect 89 511 93 523
rect 85 507 107 511
rect 97 494 101 507
rect 97 490 199 494
rect 195 486 199 490
rect 36 479 45 483
rect 167 479 174 483
rect 195 482 265 486
rect 273 482 277 496
rect 322 486 330 490
rect 424 486 432 490
rect -2 475 28 479
rect -209 457 28 461
rect 37 457 41 479
rect 273 478 282 482
rect 85 471 93 475
rect 89 465 93 471
rect 85 461 93 465
rect 101 471 107 475
rect 192 474 265 478
rect 101 465 105 471
rect 101 461 107 465
rect 36 453 45 457
rect 13 449 28 453
rect -546 324 -542 350
rect -704 320 -696 324
rect -642 320 -542 324
rect -842 284 -838 316
rect -753 312 -744 316
rect -767 308 -761 312
rect -871 283 -849 284
rect -842 283 -837 284
rect -871 282 -837 283
rect -779 282 -771 286
rect -871 280 -836 282
rect -871 -100 -867 280
rect -859 278 -836 280
rect -842 277 -837 278
rect -828 274 -819 278
rect -842 272 -836 274
rect -857 270 -836 272
rect -857 267 -837 270
rect -857 -92 -852 267
rect -841 240 -837 267
rect -828 263 -824 274
rect -775 270 -771 282
rect -766 270 -762 308
rect -753 297 -749 312
rect -700 308 -696 320
rect -704 304 -682 308
rect -693 288 -689 304
rect -546 292 -542 320
rect -717 282 -709 286
rect -693 284 -670 288
rect -662 284 -658 292
rect -612 288 -604 292
rect -550 288 -542 292
rect -713 272 -709 282
rect -662 280 -652 284
rect -693 276 -670 280
rect -779 266 -757 270
rect -770 265 -762 266
rect -770 248 -766 265
rect -770 244 -764 248
rect -756 244 -752 258
rect -707 248 -699 252
rect -756 240 -747 244
rect -841 236 -764 240
rect -756 188 -752 240
rect -703 236 -699 248
rect -693 236 -689 276
rect -662 263 -658 280
rect -608 276 -604 288
rect -612 272 -590 276
rect -600 265 -596 272
rect -645 248 -641 252
rect -546 252 -542 288
rect -636 248 -542 252
rect -707 232 -685 236
rect -546 205 -542 248
rect -231 245 -227 441
rect 0 414 28 418
rect 37 414 41 453
rect 89 449 93 461
rect 85 445 107 449
rect 99 441 103 445
rect 192 441 196 474
rect 99 437 196 441
rect 206 456 265 460
rect 273 456 277 478
rect 326 474 330 486
rect 322 470 331 474
rect 338 470 344 474
rect 326 464 330 470
rect 322 460 330 464
rect 338 464 342 470
rect 338 460 344 464
rect 85 418 93 422
rect 147 418 155 422
rect 36 410 45 414
rect -13 406 28 410
rect 37 377 41 410
rect 89 406 93 418
rect 85 402 107 406
rect 96 398 100 402
rect 206 398 210 456
rect 273 452 282 456
rect 227 448 265 452
rect 96 394 210 398
rect 273 377 277 452
rect 326 448 330 460
rect 322 444 344 448
rect 331 396 335 444
rect 546 396 551 546
rect 799 545 804 546
rect 813 542 822 546
rect 799 540 805 542
rect 784 538 805 540
rect 784 535 804 538
rect 800 508 804 535
rect 813 531 817 542
rect 866 538 870 550
rect 875 538 879 576
rect 888 565 892 580
rect 941 576 945 588
rect 937 572 959 576
rect 948 556 952 572
rect 1095 560 1099 588
rect 924 550 932 554
rect 948 552 971 556
rect 979 552 983 560
rect 1029 556 1037 560
rect 1091 556 1099 560
rect 928 540 932 550
rect 979 548 989 552
rect 948 544 971 548
rect 862 534 884 538
rect 871 533 879 534
rect 871 516 875 533
rect 871 512 877 516
rect 885 512 889 526
rect 934 516 942 520
rect 885 508 894 512
rect 800 504 877 508
rect 885 458 889 508
rect 938 504 942 516
rect 948 504 952 544
rect 979 531 983 548
rect 1033 544 1037 556
rect 1029 540 1051 544
rect 1041 533 1045 540
rect 996 516 1000 520
rect 1095 520 1099 556
rect 1005 516 1099 520
rect 934 500 956 504
rect 1095 479 1099 516
rect 884 453 889 458
rect 1091 473 1099 479
rect 1091 465 1095 473
rect 1091 453 1096 465
rect 795 429 876 433
rect 884 429 888 453
rect 1091 437 1095 453
rect 933 433 941 437
rect 995 433 1095 437
rect 795 397 799 429
rect 884 425 893 429
rect 870 421 876 425
rect 795 396 800 397
rect 331 392 551 396
rect 529 391 551 392
rect 561 395 800 396
rect 858 395 866 399
rect 561 391 801 395
rect 37 373 277 377
rect 37 267 41 373
rect 36 263 45 267
rect 167 263 174 267
rect -209 259 28 263
rect -231 241 28 245
rect 37 241 41 263
rect 85 255 93 259
rect 89 249 93 255
rect 85 245 93 249
rect 101 255 107 259
rect 101 249 105 255
rect 101 245 107 249
rect -231 52 -227 241
rect 9 233 11 237
rect 36 237 45 241
rect 16 233 28 237
rect -215 191 -214 195
rect -209 191 28 195
rect 37 191 41 237
rect 89 233 93 245
rect 237 236 241 248
rect 85 229 107 233
rect 237 232 247 236
rect 369 232 376 236
rect 97 221 101 229
rect 193 228 230 232
rect 193 221 197 228
rect 97 217 197 221
rect 205 210 230 214
rect 237 210 241 232
rect 287 224 295 228
rect 291 218 295 224
rect 287 214 295 218
rect 303 224 309 228
rect 303 218 307 224
rect 303 214 309 218
rect 85 195 93 199
rect 147 195 155 199
rect 36 187 45 191
rect -2 183 28 187
rect 37 158 41 187
rect 89 183 93 195
rect 85 179 107 183
rect 98 174 102 179
rect 205 174 209 210
rect 237 206 247 210
rect 219 202 230 206
rect 98 170 209 174
rect 237 158 241 206
rect 291 202 295 214
rect 287 198 309 202
rect 299 176 303 198
rect 299 175 411 176
rect 561 175 566 391
rect 795 390 800 391
rect 809 387 818 391
rect 795 385 801 387
rect 780 383 801 385
rect 780 380 800 383
rect 796 353 800 380
rect 809 376 813 387
rect 862 383 866 395
rect 871 383 875 421
rect 884 410 888 425
rect 937 421 941 433
rect 933 417 955 421
rect 944 401 948 417
rect 1091 405 1095 433
rect 920 395 928 399
rect 944 397 967 401
rect 975 397 979 405
rect 1025 401 1033 405
rect 1087 401 1095 405
rect 924 385 928 395
rect 975 393 985 397
rect 944 389 967 393
rect 858 379 880 383
rect 867 378 875 379
rect 867 361 871 378
rect 867 357 873 361
rect 881 357 885 371
rect 930 361 938 365
rect 881 353 890 357
rect 796 349 873 353
rect 792 271 873 275
rect 881 271 885 353
rect 934 349 938 361
rect 944 349 948 389
rect 975 376 979 393
rect 1029 389 1033 401
rect 1025 385 1047 389
rect 1037 378 1041 385
rect 992 361 996 365
rect 1091 365 1095 401
rect 1001 361 1095 365
rect 930 345 952 349
rect 1091 324 1095 361
rect 1088 318 1095 324
rect 1088 279 1092 318
rect 930 275 938 279
rect 992 275 1092 279
rect 792 239 796 271
rect 881 267 890 271
rect 867 263 873 267
rect 792 238 797 239
rect 299 172 566 175
rect 400 170 566 172
rect 575 237 797 238
rect 855 237 863 241
rect 575 233 798 237
rect 37 154 241 158
rect -231 48 29 52
rect 37 48 41 154
rect 86 52 94 56
rect 148 52 156 56
rect 37 44 46 48
rect 15 40 29 44
rect 37 30 41 44
rect 90 40 94 52
rect 86 36 108 40
rect 99 33 103 36
rect 260 33 268 37
rect 322 33 330 37
rect 99 29 203 33
rect 211 25 220 29
rect 202 21 203 25
rect 264 21 268 33
rect 260 17 282 21
rect 271 4 275 17
rect 271 3 389 4
rect 575 3 580 233
rect 792 232 797 233
rect 806 229 815 233
rect 792 227 798 229
rect 777 225 798 227
rect 777 222 797 225
rect 793 195 797 222
rect 806 218 810 229
rect 859 225 863 237
rect 868 225 872 263
rect 881 252 885 267
rect 934 263 938 275
rect 930 259 952 263
rect 941 243 945 259
rect 1088 247 1092 275
rect 917 237 925 241
rect 941 239 964 243
rect 972 239 976 247
rect 1022 243 1030 247
rect 1084 243 1092 247
rect 921 227 925 237
rect 972 235 982 239
rect 941 231 964 235
rect 855 221 877 225
rect 864 220 872 221
rect 864 203 868 220
rect 864 199 870 203
rect 878 199 882 213
rect 927 203 935 207
rect 878 195 887 199
rect 793 191 870 195
rect 789 67 870 71
rect 878 67 882 195
rect 931 191 935 203
rect 941 191 945 231
rect 972 218 976 235
rect 1026 231 1030 243
rect 1022 227 1044 231
rect 1034 220 1038 227
rect 989 203 993 207
rect 1088 207 1092 243
rect 998 203 1092 207
rect 927 187 949 191
rect 1088 106 1092 203
rect 1084 102 1092 106
rect 1085 101 1092 102
rect 1085 75 1089 101
rect 927 71 935 75
rect 989 71 1089 75
rect 789 35 793 67
rect 878 63 887 67
rect 864 59 870 63
rect 789 34 794 35
rect 772 33 794 34
rect 852 33 860 37
rect 772 29 795 33
rect 789 28 794 29
rect 803 25 812 29
rect 789 23 795 25
rect 774 21 795 23
rect 774 18 794 21
rect 271 0 580 3
rect 379 -2 580 0
rect 790 -9 794 18
rect 803 14 807 25
rect 856 21 860 33
rect 865 21 869 59
rect 878 48 882 63
rect 931 59 935 71
rect 927 55 949 59
rect 938 39 942 55
rect 1085 43 1089 71
rect 914 33 922 37
rect 938 35 961 39
rect 969 35 973 43
rect 1019 39 1027 43
rect 1081 39 1089 43
rect 918 23 922 33
rect 969 31 979 35
rect 938 27 961 31
rect 852 17 874 21
rect 861 16 869 17
rect 861 -1 865 16
rect 861 -5 867 -1
rect 875 -5 879 9
rect 924 -1 932 3
rect 875 -9 884 -5
rect 790 -13 867 -9
rect 875 -61 879 -9
rect 928 -13 932 -1
rect 938 -13 942 27
rect 969 14 973 31
rect 1023 27 1027 39
rect 1019 23 1041 27
rect 1031 16 1035 23
rect 986 -1 990 3
rect 1085 3 1089 39
rect 995 -1 1089 3
rect 924 -17 946 -13
rect 1085 -44 1089 -1
rect -633 -92 -625 -88
rect -571 -92 -563 -88
rect -857 -96 -690 -92
rect -857 -97 -691 -96
rect -682 -100 -673 -96
rect -871 -104 -690 -100
rect -629 -104 -625 -92
rect -633 -108 -611 -104
rect -622 -141 -618 -108
rect -622 -145 -39 -141
<< m2contact >>
rect -168 1304 -163 1310
rect -159 1215 -154 1221
rect -128 1106 -123 1112
rect 295 1007 300 1012
rect -740 965 -735 970
rect -650 965 -645 970
rect -700 940 -695 945
rect -815 931 -810 936
rect -743 931 -738 936
rect -650 931 -645 936
rect -587 933 -582 938
rect -628 921 -623 926
rect 0 927 5 932
rect 6 909 11 914
rect 279 924 284 929
rect -214 901 -209 906
rect -743 809 -738 814
rect -653 809 -648 814
rect -703 784 -698 789
rect -818 775 -813 780
rect -746 775 -741 780
rect -653 775 -648 780
rect -590 777 -585 782
rect -631 765 -626 770
rect -747 654 -742 659
rect -657 654 -652 659
rect -707 629 -702 634
rect -822 620 -817 625
rect -750 620 -745 625
rect -657 620 -652 625
rect -594 622 -589 627
rect -635 610 -630 615
rect -750 496 -745 501
rect -660 496 -655 501
rect -710 471 -705 476
rect -825 462 -820 467
rect -753 462 -748 467
rect -660 462 -655 467
rect -597 464 -592 469
rect -638 452 -633 457
rect 10 875 15 880
rect -7 821 -2 826
rect 3 813 8 818
rect 10 786 15 791
rect -2 751 3 756
rect 1 733 6 738
rect 10 725 15 730
rect 6 690 11 695
rect 295 754 300 759
rect 891 716 896 721
rect 981 716 986 721
rect 931 691 936 696
rect 816 682 821 687
rect 888 682 893 687
rect 269 642 274 647
rect -13 545 -8 550
rect 981 682 986 687
rect 1044 684 1049 689
rect 1003 672 1008 677
rect -214 537 -209 542
rect 7 511 12 516
rect -7 475 -2 480
rect -214 456 -209 461
rect 8 449 13 454
rect -231 441 -226 446
rect -753 292 -748 297
rect -663 292 -658 297
rect -713 267 -708 272
rect -828 258 -823 263
rect -756 258 -751 263
rect -663 258 -658 263
rect -600 260 -595 265
rect -641 248 -636 253
rect -5 414 0 419
rect -18 405 -13 410
rect 222 447 227 452
rect 888 560 893 565
rect 978 560 983 565
rect 928 535 933 540
rect 813 526 818 531
rect 885 526 890 531
rect 978 526 983 531
rect 1041 528 1046 533
rect 1000 516 1005 521
rect -214 259 -209 264
rect 11 233 16 238
rect -214 191 -209 196
rect -7 183 -2 188
rect 214 201 219 206
rect 884 405 889 410
rect 974 405 979 410
rect 924 380 929 385
rect 809 371 814 376
rect 881 371 886 376
rect 974 371 979 376
rect 1037 373 1042 378
rect 996 361 1001 366
rect 10 40 15 45
rect 197 21 202 26
rect 881 247 886 252
rect 971 247 976 252
rect 921 222 926 227
rect 806 213 811 218
rect 878 213 883 218
rect 971 213 976 218
rect 1034 215 1039 220
rect 993 203 998 208
rect 878 43 883 48
rect 968 43 973 48
rect 918 18 923 23
rect 803 9 808 14
rect 875 9 880 14
rect 968 9 973 14
rect 1031 11 1036 16
rect 990 -1 995 4
<< metal2 >>
rect -169 1304 -168 1308
rect -167 1287 -163 1304
rect -159 1172 -155 1215
rect -159 1164 -155 1167
rect -128 1099 -124 1106
rect 300 1007 342 1011
rect -735 965 -650 970
rect -695 940 -625 943
rect -810 931 -743 936
rect -738 931 -650 936
rect -628 926 -625 940
rect -587 914 -583 933
rect -174 927 0 931
rect -587 910 -512 914
rect -192 909 6 913
rect -738 809 -653 814
rect -698 784 -628 787
rect -813 775 -746 780
rect -741 775 -653 780
rect -631 770 -628 784
rect -590 758 -586 777
rect -515 758 -490 759
rect -590 754 -490 758
rect -742 654 -657 659
rect -702 629 -632 632
rect -817 620 -750 625
rect -745 620 -657 625
rect -635 615 -632 629
rect -594 603 -590 622
rect -519 603 -514 604
rect -214 603 -210 901
rect 279 896 283 924
rect 269 892 283 896
rect -162 875 10 879
rect -174 821 -7 825
rect -192 813 3 817
rect -153 787 10 791
rect -174 751 -2 755
rect -192 733 1 737
rect -123 725 10 729
rect -174 690 6 694
rect 269 647 273 892
rect 338 881 342 1007
rect 279 877 342 881
rect 279 759 283 877
rect 279 755 295 759
rect 294 754 295 755
rect 896 716 981 721
rect 936 691 1006 694
rect 821 682 888 687
rect 893 682 981 687
rect 1003 677 1006 691
rect 1044 665 1048 684
rect 1119 665 1124 666
rect 1044 661 1124 665
rect -594 599 -210 603
rect -214 542 -210 599
rect -192 545 -13 549
rect -745 496 -660 501
rect -705 471 -635 474
rect -820 462 -753 467
rect -748 462 -660 467
rect -638 457 -635 471
rect -597 445 -593 464
rect -214 461 -210 537
rect -162 511 7 515
rect -192 475 -7 479
rect -522 445 -517 446
rect -597 441 -231 445
rect -748 292 -663 297
rect -708 267 -638 270
rect -823 258 -756 263
rect -751 258 -663 263
rect -641 253 -638 267
rect -214 264 -210 456
rect -153 449 8 453
rect 223 452 227 627
rect 893 560 978 565
rect 933 535 1003 538
rect 818 526 885 531
rect 890 526 978 531
rect 1000 521 1003 535
rect 1041 509 1045 528
rect 1116 509 1121 510
rect 1041 505 1121 509
rect 221 447 222 451
rect -192 414 -5 418
rect -123 406 -18 410
rect -29 400 -25 406
rect 889 405 974 410
rect 929 380 999 383
rect 814 371 881 376
rect 886 371 974 376
rect 996 366 999 380
rect 1037 354 1041 373
rect 1112 354 1117 355
rect 1037 350 1117 354
rect -600 241 -596 260
rect -525 241 -520 242
rect -600 237 -520 241
rect -214 196 -210 259
rect -162 233 11 237
rect 214 206 218 307
rect 886 247 971 252
rect 926 222 996 225
rect 811 213 878 218
rect 883 213 971 218
rect 993 208 996 222
rect 213 201 214 205
rect 1034 196 1038 215
rect 1109 196 1114 197
rect 1034 192 1114 196
rect -214 190 -210 191
rect -153 183 -7 187
rect -17 177 -13 183
rect -163 40 10 44
rect 197 26 201 84
rect 883 43 968 48
rect 923 18 993 21
rect 808 9 875 14
rect 880 9 968 14
rect 990 4 993 18
rect 1031 -8 1035 11
rect 1106 -8 1111 -7
rect 1031 -12 1111 -8
<< m3contact >>
rect -167 1282 -162 1287
rect -159 1167 -154 1172
rect -128 1094 -123 1099
rect -179 927 -174 932
rect -512 910 -507 915
rect -197 909 -192 914
rect -490 754 -485 759
rect -167 875 -162 880
rect -179 821 -174 826
rect -197 813 -192 818
rect -158 786 -153 791
rect -179 751 -174 756
rect -197 733 -192 738
rect -128 724 -123 729
rect -179 690 -174 695
rect -197 545 -192 550
rect -167 511 -162 516
rect -197 475 -192 480
rect -158 449 -153 454
rect -197 414 -192 419
rect -128 405 -123 410
rect -167 233 -162 238
rect -158 183 -153 188
rect -168 40 -163 45
<< metal3 >>
rect -260 948 -174 953
rect -513 915 -506 916
rect -260 915 -255 948
rect -179 932 -174 948
rect -513 910 -512 915
rect -507 910 -255 915
rect -197 914 -192 919
rect -513 909 -506 910
rect -197 818 -192 909
rect -491 759 -484 760
rect -197 759 -192 813
rect -491 754 -490 759
rect -485 754 -192 759
rect -491 753 -484 754
rect -197 738 -192 754
rect -197 550 -192 733
rect -179 826 -174 927
rect -179 756 -174 821
rect -179 695 -174 751
rect -167 880 -164 1282
rect -197 480 -192 545
rect -197 419 -192 475
rect -197 197 -192 414
rect -167 516 -164 875
rect -158 791 -155 1167
rect -128 1093 -123 1094
rect -167 238 -164 511
rect -158 454 -155 786
rect -128 729 -125 1093
rect -167 45 -164 233
rect -158 188 -155 449
rect -128 410 -125 724
rect -128 399 -125 405
rect -158 178 -155 183
rect -167 14 -164 40
<< labels >>
rlabel metal1 384 0 388 4 1 c2
rlabel metal1 405 172 409 176 1 c3
rlabel metal1 518 392 522 396 1 c4
rlabel metal1 562 705 566 709 1 c5
rlabel metal1 -756 188 -752 192 1 vdd
rlabel metal1 -546 205 -542 209 1 gnd
rlabel metal1 -859 278 -854 283 3 a0
rlabel metal1 -857 267 -852 272 3 b0
rlabel metal1 -854 471 -849 476 1 b1
rlabel metal1 -856 482 -851 487 1 a1
rlabel metal1 -851 629 -846 634 1 b2
rlabel metal1 -853 640 -848 645 1 a2
rlabel metal1 -847 784 -842 789 1 b3
rlabel metal1 -849 795 -844 800 1 a3
rlabel metal1 -844 940 -839 945 1 b4
rlabel metal1 -846 951 -841 956 1 a4
rlabel metal1 -567 -92 -563 -88 7 gnd
rlabel metal1 -682 -100 -678 -96 7 vdd
rlabel metal1 -696 -96 -692 -92 3 b
rlabel metal1 -696 -104 -692 -100 3 a
rlabel metal1 -622 -108 -618 -104 7 out
rlabel metal1 218 1046 222 1050 7 vdd
rlabel metal1 204 1050 208 1054 3 b
rlabel metal1 204 1042 208 1046 3 a
rlabel metal1 333 1054 337 1058 7 gnd
rlabel metal1 278 1038 282 1042 7 out
rlabel metal1 306 755 309 759 1 g4
rlabel m2contact 10 725 13 729 1 g2
rlabel m2contact 10 875 13 879 1 g0
rlabel m2contact 10 787 13 791 1 g1
rlabel metal1 10 511 13 515 1 g0
rlabel metal1 10 519 13 523 1 p1
rlabel metal1 10 537 13 541 1 p2
rlabel metal1 10 545 13 549 1 p3
rlabel metal1 10 733 13 737 1 p3
rlabel metal1 10 795 13 799 1 p2
rlabel metal1 10 901 13 905 1 p2
rlabel metal1 10 883 13 887 1 p1
rlabel metal1 10 909 13 913 1 p3
rlabel metal1 10 927 13 931 1 p4
rlabel metal1 10 259 13 263 1 p2
rlabel metal1 24 241 27 245 1 p1
rlabel metal1 24 233 27 237 1 g0
rlabel metal1 24 821 27 825 1 p4
rlabel metal1 24 813 27 817 1 p3
rlabel metal1 24 751 27 755 1 p4
rlabel metal1 24 690 27 694 1 p4
rlabel metal1 24 475 27 479 1 p3
rlabel metal1 24 457 27 461 1 p2
rlabel metal1 24 414 27 418 1 p3
rlabel metal1 24 191 27 195 1 p2
rlabel metal1 24 48 27 52 1 p1
rlabel metal1 24 183 27 187 1 g1
rlabel metal1 24 406 27 410 1 g2
rlabel metal1 24 449 27 453 1 g1
rlabel metal1 24 682 27 686 1 g3
rlabel metal1 24 40 27 44 1 g0
rlabel metal1 260 448 263 452 1 g3
rlabel metal1 225 202 228 206 1 g2
rlabel m2contact 197 21 200 25 1 g1
rlabel metal1 875 -61 879 -57 1 vdd
rlabel metal1 1085 -44 1089 -40 1 gnd
rlabel metal2 1106 -12 1111 -7 1 p0
rlabel metal1 772 29 777 34 3 a0
rlabel metal1 774 18 779 23 3 b0
rlabel metal1 777 222 782 227 1 b1
rlabel metal1 775 233 780 238 1 a1
rlabel metal1 780 380 785 385 1 b2
rlabel metal1 778 391 783 396 1 a2
rlabel metal1 784 535 789 540 1 b3
rlabel metal1 782 546 787 551 1 a3
rlabel metal1 787 691 792 696 1 b4
rlabel metal1 785 702 790 707 1 a4
rlabel metal2 1119 661 1124 666 7 p4
rlabel metal2 1116 505 1121 510 1 p3
rlabel metal2 1112 350 1117 355 1 p2
rlabel metal2 1109 192 1114 197 1 p1
rlabel metal1 -189 1154 -185 1158 7 vdd
rlabel metal1 -203 1158 -199 1162 3 b
rlabel metal1 -203 1150 -199 1154 3 a
rlabel metal1 -74 1162 -70 1166 7 gnd
rlabel metal1 -129 1146 -125 1150 7 out
rlabel metal1 -159 1270 -155 1274 7 out
rlabel metal1 -104 1286 -100 1290 7 gnd
rlabel metal1 -233 1274 -229 1278 3 a
rlabel metal1 -233 1282 -229 1286 3 b
rlabel metal1 -219 1278 -215 1282 7 vdd
rlabel metal1 -169 1405 -165 1409 7 out
rlabel metal1 -229 1413 -225 1417 7 vdd
rlabel metal1 -114 1421 -110 1425 7 gnd
rlabel metal1 -243 1409 -239 1413 3 a
rlabel metal1 -243 1417 -239 1421 3 b
<< end >>
