magic
tech scmos
timestamp 1763386966
<< nwell >>
rect -11 71 52 123
<< ntransistor >>
rect 0 -25 2 55
rect 8 -25 10 55
rect 31 -25 33 55
rect 39 -25 41 55
<< ptransistor >>
rect 0 77 2 117
rect 8 77 10 117
rect 31 77 33 117
rect 39 77 41 117
<< ndiffusion >>
rect -1 -25 0 55
rect 2 -25 3 55
rect 7 -25 8 55
rect 10 -25 11 55
rect 30 -25 31 55
rect 33 -25 34 55
rect 38 -25 39 55
rect 41 -25 42 55
<< pdiffusion >>
rect -1 77 0 117
rect 2 77 3 117
rect 7 77 8 117
rect 10 77 11 117
rect 30 77 31 117
rect 33 77 34 117
rect 38 77 39 117
rect 41 77 42 117
<< ndcontact >>
rect -5 -25 -1 55
rect 3 -25 7 55
rect 11 -25 15 55
rect 26 -25 30 55
rect 34 -25 38 55
rect 42 -25 46 55
<< pdcontact >>
rect -5 77 -1 117
rect 3 77 7 117
rect 11 77 15 117
rect 26 77 30 117
rect 34 77 38 117
rect 42 77 46 117
<< polysilicon >>
rect 0 117 2 130
rect 8 117 10 130
rect 31 117 33 130
rect 39 117 41 130
rect 0 55 2 77
rect 8 55 10 77
rect 31 55 33 77
rect 39 55 41 77
rect 0 -30 2 -25
rect 8 -30 10 -25
rect 31 -30 33 -25
rect 39 -30 41 -25
<< polycontact >>
rect -1 130 3 134
rect 7 130 11 134
rect 30 130 34 134
rect 38 130 42 134
<< metal1 >>
rect -1 134 3 140
rect 7 134 11 140
rect 30 134 34 140
rect 38 134 42 140
rect 3 117 7 126
rect 34 117 38 126
rect -5 73 -1 77
rect 11 73 15 77
rect 26 73 30 77
rect 42 73 46 77
rect -5 69 16 73
rect 21 69 46 73
rect -5 55 -1 69
rect 26 68 30 69
rect 11 57 16 61
rect 21 57 30 61
rect 11 55 15 57
rect 26 55 30 57
rect 42 -33 46 -25
<< labels >>
rlabel metal1 3 122 7 126 1 vdd
rlabel metal1 7 136 11 140 5 b
rlabel metal1 -1 136 3 140 5 a
rlabel metal1 -5 62 -1 66 1 out
rlabel metal1 42 -33 46 -29 1 gnd
rlabel metal1 30 136 34 140 5 a
rlabel metal1 38 136 42 140 5 b
rlabel metal1 34 122 38 126 1 vdd
<< end >>
