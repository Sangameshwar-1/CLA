* Test file for 4-input NAND gate (Magic extracted)
* ==========================================================

.include "/home/sangam/Documents/VLSI_PROJ_2017/MAGIC/TSMC_180nm.txt"

* SPICE3 file created from nand_4.ext - technology: scmos
.option scale=0.09u

.subckt nand4 a b c d out vdd Gnd

* SPICE3 file created from nand_4.ext - technology: scmos

.option scale=0.09u

M1000 out d vdd w_n11_71# CMOSP w=40 l=2
+  ad=800 pd=360 as=480 ps=184
M1001 gnd d a_28_n25# Gnd CMOSN w=80 l=2
+  ad=400 pd=170 as=480 ps=172
M1002 a_10_n25# b a_2_n25# Gnd CMOSN w=80 l=2
+  ad=800 pd=340 as=480 ps=172
M1003 vdd a out w_n11_71# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_2_n25# a out Gnd CMOSN w=80 l=2
+  ad=0 pd=0 as=400 ps=170
M1005 vdd c out w_n11_71# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 out b vdd w_n11_71# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 a_28_n25# c a_10_n25# Gnd CMOSN w=80 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vdd w_n11_71# 0.07fF
C1 b a 0.27fF
C2 a_28_n25# a_10_n25# 0.82fF
C3 d c 0.27fF
C4 a out 0.08fF
C5 d out 0.08fF
C6 b out 0.08fF
C7 c out 0.08fF
C8 a_10_n25# a_2_n25# 0.82fF
C9 a_2_n25# out 0.82fF
C10 a_10_n25# out 0.02fF
C11 b vdd 0.10fF
C12 vdd c 0.10fF
C13 vdd out 1.79fF
C14 a_28_n25# gnd 0.82fF
C15 w_n11_71# a 0.08fF
C16 d w_n11_71# 0.08fF
C17 b w_n11_71# 0.08fF
C18 w_n11_71# c 0.08fF
C19 w_n11_71# out 0.28fF
C20 gnd Gnd 0.11fF
C21 a_28_n25# Gnd 0.01fF
C22 a_10_n25# Gnd 0.23fF
C23 a_2_n25# Gnd 0.01fF
C24 vdd Gnd 0.06fF
C25 out Gnd 0.12fF
C26 d Gnd 0.12fF
C27 c Gnd 0.12fF
C28 b Gnd 0.12fF
C29 a Gnd 0.12fF
C30 w_n11_71# Gnd 3.03fF



.ends nand4

* ========== TESTBENCH ==========

.param SUPPLY=1.8
.global gnd vdd

VDD vdd gnd {SUPPLY}

* Truth Table for 4-input NAND
* A B C D | OUT
* 0 0 0 0 | 1
* 0 0 0 1 | 1
* ... (14 more combinations)
* 1 1 1 1 | 0

* Test 1: A=0, B=0, C=0, D=0 -> OUT=1
VA_0000 a_0000 gnd 0
VB_0000 b_0000 gnd 0
VC_0000 c_0000 gnd 0
VD_0000 d_0000 gnd 0
Xnand_0000 a_0000 b_0000 c_0000 d_0000 out_0000 vdd gnd nand4
Cload_0000 out_0000 gnd 10f

* Test 2: A=0, B=0, C=0, D=1 -> OUT=1
VA_0001 a_0001 gnd 0
VB_0001 b_0001 gnd 0
VC_0001 c_0001 gnd 0
VD_0001 d_0001 gnd {SUPPLY}
Xnand_0001 a_0001 b_0001 c_0001 d_0001 out_0001 vdd gnd nand4
Cload_0001 out_0001 gnd 10f

* Test 3: A=0, B=1, C=1, D=1 -> OUT=1
VA_0111 a_0111 gnd 0
VB_0111 b_0111 gnd {SUPPLY}
VC_0111 c_0111 gnd {SUPPLY}
VD_0111 d_0111 gnd {SUPPLY}
Xnand_0111 a_0111 b_0111 c_0111 d_0111 out_0111 vdd gnd nand4
Cload_0111 out_0111 gnd 10f

* Test 4: A=1, B=0, C=1, D=1 -> OUT=1
VA_1011 a_1011 gnd {SUPPLY}
VB_1011 b_1011 gnd 0
VC_1011 c_1011 gnd {SUPPLY}
VD_1011 d_1011 gnd {SUPPLY}
Xnand_1011 a_1011 b_1011 c_1011 d_1011 out_1011 vdd gnd nand4
Cload_1011 out_1011 gnd 10f

* Test 5: A=1, B=1, C=0, D=1 -> OUT=1
VA_1101 a_1101 gnd {SUPPLY}
VB_1101 b_1101 gnd {SUPPLY}
VC_1101 c_1101 gnd 0
VD_1101 d_1101 gnd {SUPPLY}
Xnand_1101 a_1101 b_1101 c_1101 d_1101 out_1101 vdd gnd nand4
Cload_1101 out_1101 gnd 10f

* Test 6: A=1, B=1, C=1, D=0 -> OUT=1
VA_1110 a_1110 gnd {SUPPLY}
VB_1110 b_1110 gnd {SUPPLY}
VC_1110 c_1110 gnd {SUPPLY}
VD_1110 d_1110 gnd 0
Xnand_1110 a_1110 b_1110 c_1110 d_1110 out_1110 vdd gnd nand4
Cload_1110 out_1110 gnd 10f

* Test 7: A=1, B=1, C=1, D=1 -> OUT=0
VA_1111 a_1111 gnd {SUPPLY}
VB_1111 b_1111 gnd {SUPPLY}
VC_1111 c_1111 gnd {SUPPLY}
VD_1111 d_1111 gnd {SUPPLY}
Xnand_1111 a_1111 b_1111 c_1111 d_1111 out_1111 vdd gnd nand4
Cload_1111 out_1111 gnd 10f

* Dynamic test with pulses
VA_dyn a_dyn gnd PULSE(0 {SUPPLY} 1n 100p 100p 4n 8n)
VB_dyn b_dyn gnd PULSE(0 {SUPPLY} 2n 100p 100p 8n 16n)
VC_dyn c_dyn gnd PULSE(0 {SUPPLY} 4n 100p 100p 16n 32n)
VD_dyn d_dyn gnd PULSE(0 {SUPPLY} 8n 100p 100p 32n 64n)
Xnand_dyn a_dyn b_dyn c_dyn d_dyn out_dyn vdd gnd nand4
Cload_dyn out_dyn gnd 10f

.control
set numdgt=12

echo ""
echo "=========================================="
echo "  4-INPUT NAND GATE TRUTH TABLE TEST"
echo "=========================================="
echo "  (Magic Extracted Layout with TSMC 180nm)"
echo ""

* DC Operating Point
op

echo "Truth Table Verification (selected cases):"
echo "  A B C D | OUT | Expected"
echo "  --------+-----+---------"

* Test 0000
let v_0000 = v(out_0000)
if v_0000 > 1.5
    echo "  0 0 0 0 |  1  |    1     PASS"
else
    echo "  0 0 0 0 |  0  |    1     FAIL"
end

* Test 0001
let v_0001 = v(out_0001)
if v_0001 > 1.5
    echo "  0 0 0 1 |  1  |    1     PASS"
else
    echo "  0 0 0 1 |  0  |    1     FAIL"
end

* Test 0111
let v_0111 = v(out_0111)
if v_0111 > 1.5
    echo "  0 1 1 1 |  1  |    1     PASS"
else
    echo "  0 1 1 1 |  0  |    1     FAIL"
end

* Test 1011
let v_1011 = v(out_1011)
if v_1011 > 1.5
    echo "  1 0 1 1 |  1  |    1     PASS"
else
    echo "  1 0 1 1 |  0  |    1     FAIL"
end

* Test 1101
let v_1101 = v(out_1101)
if v_1101 > 1.5
    echo "  1 1 0 1 |  1  |    1     PASS"
else
    echo "  1 1 0 1 |  0  |    1     FAIL"
end

* Test 1110
let v_1110 = v(out_1110)
if v_1110 > 1.5
    echo "  1 1 1 0 |  1  |    1     PASS"
else
    echo "  1 1 1 0 |  0  |    1     FAIL"
end

* Test 1111
let v_1111 = v(out_1111)
if v_1111 < 0.3
    echo "  1 1 1 1 |  0  |    0     PASS"
else
    echo "  1 1 1 1 |  1  |    0     FAIL"
end

echo ""
echo "=========================================="
echo "  DYNAMIC TRANSIENT ANALYSIS"
echo "=========================================="
echo ""

tran 10p 40n

* Measure propagation delays (worst case: all inputs high -> low)
meas tran tpHL TRIG v(a_dyn) VAL=0.9 RISE=1 TARG v(out_dyn) VAL=0.9 FALL=1
meas tran tpLH TRIG v(a_dyn) VAL=0.9 FALL=1 TARG v(out_dyn) VAL=0.9 RISE=1
let tpd_avg = (tpHL + tpLH) / 2

echo "Timing Characteristics:"
echo "  tpHL (High->Low): " $&tpHL "s"
echo "  tpLH (Low->High): " $&tpLH "s"
echo "  tpd (Average):    " $&tpd_avg "s"
echo ""

* Rise and fall times
meas tran tr TRIG v(out_dyn) VAL=0.18 RISE=1 TARG v(out_dyn) VAL=1.62 RISE=1
meas tran tf TRIG v(out_dyn) VAL=1.62 FALL=1 TARG v(out_dyn) VAL=0.18 FALL=1

echo "Edge Rates:"
echo "  Rise time (10%-90%): " $&tr "s"
echo "  Fall time (90%-10%): " $&tf "s"
echo ""

* Measure power
meas tran iavg AVG i(VDD) FROM=2n TO=40n
let pavg = abs(iavg) * 1.8
echo "Power Consumption:"
echo "  Average Power: " $&pavg "W"
echo ""

echo "=========================================="
echo "  Layout Extracted - Includes Parasitics"
echo "=========================================="
echo ""

* Plot waveforms
plot v(a_dyn) v(b_dyn)+2 v(c_dyn)+4 v(d_dyn)+6 v(out_dyn)+8

* Detailed view of first transition
plot v(a_dyn) v(b_dyn)+2 v(c_dyn)+4 v(d_dyn)+6 v(out_dyn)+8 xlimit 0 10n

.endc
.end
