magic
tech scmos
timestamp 1763547437
<< nwell >>
rect 682 681 734 713
rect 774 679 826 681
rect 607 643 659 675
rect 773 647 826 679
rect 679 609 731 641
<< ntransistor >>
rect 750 700 790 702
rect 750 692 790 694
rect 842 668 882 670
rect 675 662 715 664
rect 842 660 882 662
rect 675 654 715 656
rect 747 628 787 630
rect 747 620 787 622
<< ptransistor >>
rect 688 700 728 702
rect 688 692 728 694
rect 780 668 820 670
rect 613 662 653 664
rect 780 660 820 662
rect 613 654 653 656
rect 685 628 725 630
rect 685 620 725 622
<< ndiffusion >>
rect 750 702 790 703
rect 750 699 790 700
rect 750 694 790 695
rect 750 691 790 692
rect 842 670 882 671
rect 675 664 715 665
rect 675 661 715 662
rect 842 667 882 668
rect 842 662 882 663
rect 675 656 715 657
rect 842 659 882 660
rect 675 653 715 654
rect 747 630 787 631
rect 747 627 787 628
rect 747 622 787 623
rect 747 619 787 620
<< pdiffusion >>
rect 688 702 728 703
rect 688 699 728 700
rect 688 694 728 695
rect 688 691 728 692
rect 613 664 653 665
rect 780 670 820 671
rect 780 667 820 668
rect 613 661 653 662
rect 613 656 653 657
rect 780 662 820 663
rect 780 659 820 660
rect 613 653 653 654
rect 685 630 725 631
rect 685 627 725 628
rect 685 622 725 623
rect 685 619 725 620
<< ndcontact >>
rect 750 703 790 707
rect 750 695 790 699
rect 750 687 790 691
rect 675 665 715 669
rect 842 671 882 675
rect 675 657 715 661
rect 842 663 882 667
rect 842 655 882 659
rect 675 649 715 653
rect 747 631 787 635
rect 747 623 787 627
rect 747 615 787 619
<< pdcontact >>
rect 688 703 728 707
rect 688 695 728 699
rect 688 687 728 691
rect 780 671 820 675
rect 613 665 653 669
rect 780 663 820 667
rect 613 657 653 661
rect 780 655 820 659
rect 613 649 653 653
rect 685 631 725 635
rect 685 623 725 627
rect 685 615 725 619
<< polysilicon >>
rect 675 700 688 702
rect 728 700 750 702
rect 790 700 793 702
rect 675 692 688 694
rect 728 692 750 694
rect 790 692 793 694
rect 766 668 780 670
rect 820 668 842 670
rect 882 668 885 670
rect 600 662 613 664
rect 653 662 675 664
rect 715 662 718 664
rect 766 660 780 662
rect 820 660 842 662
rect 882 660 885 662
rect 600 654 613 656
rect 653 654 675 656
rect 715 654 718 656
rect 672 628 685 630
rect 725 628 747 630
rect 787 628 790 630
rect 672 620 685 622
rect 725 620 747 622
rect 787 620 790 622
<< polycontact >>
rect 671 699 675 703
rect 671 691 675 695
rect 596 661 600 665
rect 762 667 766 671
rect 596 653 600 657
rect 762 659 766 663
rect 668 627 672 631
rect 668 619 672 623
<< metal1 >>
rect 590 699 671 703
rect 679 699 683 728
rect 886 707 890 725
rect 728 703 736 707
rect 790 703 890 707
rect 590 667 594 699
rect 679 695 688 699
rect 665 691 671 695
rect 590 666 595 667
rect 573 665 595 666
rect 653 665 661 669
rect 573 661 596 665
rect 590 660 595 661
rect 604 657 613 661
rect 590 655 596 657
rect 575 653 596 655
rect 575 650 595 653
rect 591 623 595 650
rect 604 646 608 657
rect 657 653 661 665
rect 666 653 670 691
rect 679 680 683 695
rect 732 691 736 703
rect 728 687 750 691
rect 739 671 743 687
rect 886 675 890 703
rect 715 665 723 669
rect 739 667 762 671
rect 770 667 774 675
rect 820 671 828 675
rect 882 671 890 675
rect 719 655 723 665
rect 770 663 780 667
rect 739 659 762 663
rect 653 649 675 653
rect 662 648 670 649
rect 662 631 666 648
rect 662 627 668 631
rect 676 627 680 641
rect 725 631 733 635
rect 676 623 685 627
rect 591 619 668 623
rect 676 546 680 623
rect 729 619 733 631
rect 739 619 743 659
rect 770 646 774 663
rect 824 659 828 671
rect 820 655 842 659
rect 832 648 836 655
rect 787 631 791 635
rect 886 635 890 671
rect 796 631 890 635
rect 725 615 747 619
rect 886 588 890 631
rect 676 542 681 546
<< m2contact >>
rect 679 675 684 680
rect 769 675 774 680
rect 719 650 724 655
rect 604 641 609 646
rect 676 641 681 646
rect 769 641 774 646
rect 832 643 837 648
rect 791 631 796 636
<< metal2 >>
rect 684 675 769 680
rect 724 650 794 653
rect 609 641 676 646
rect 681 641 769 646
rect 791 636 794 650
rect 832 624 836 643
rect 907 624 912 625
rect 832 620 912 624
rect 1252 579 1264 583
<< labels >>
rlabel metal1 676 579 680 583 1 vdd
rlabel metal2 907 620 911 624 7 xor
rlabel metal1 886 588 890 592 1 gnd
rlabel metal1 590 650 595 657 3 b
rlabel metal1 590 660 595 667 3 a
rlabel metal2 1259 579 1264 583 7 xorabc
<< end >>
