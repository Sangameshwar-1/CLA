magic
tech scmos
timestamp 1763552233
<< nwell >>
rect 4 993 56 1072
rect 4 905 56 963
rect 4 843 56 893
rect 286 873 338 952
rect 4 800 56 832
rect 4 629 56 687
rect 4 567 56 617
rect 241 566 293 624
rect 4 524 56 556
rect 4 351 56 401
rect 4 301 56 333
rect 206 320 258 370
rect 5 158 57 190
rect 179 139 231 171
<< ntransistor >>
rect 72 1056 172 1058
rect 72 1038 172 1040
rect 72 1030 172 1032
rect 72 1012 172 1014
rect 72 1004 172 1006
rect 72 950 152 952
rect 72 942 152 944
rect 354 936 454 938
rect 72 924 152 926
rect 72 916 152 918
rect 354 918 454 920
rect 354 910 454 912
rect 354 892 454 894
rect 354 884 454 886
rect 72 880 132 882
rect 72 862 132 864
rect 72 854 132 856
rect 72 819 112 821
rect 72 811 112 813
rect 72 674 152 676
rect 72 666 152 668
rect 72 648 152 650
rect 72 640 152 642
rect 309 611 389 613
rect 72 604 132 606
rect 309 603 389 605
rect 72 586 132 588
rect 309 585 389 587
rect 72 578 132 580
rect 309 577 389 579
rect 72 543 112 545
rect 72 535 112 537
rect 72 388 132 390
rect 72 370 132 372
rect 72 362 132 364
rect 274 357 334 359
rect 274 339 334 341
rect 274 331 334 333
rect 72 320 112 322
rect 72 312 112 314
rect 73 177 113 179
rect 73 169 113 171
rect 247 158 287 160
rect 247 150 287 152
<< ptransistor >>
rect 10 1056 50 1058
rect 10 1038 50 1040
rect 10 1030 50 1032
rect 10 1012 50 1014
rect 10 1004 50 1006
rect 10 950 50 952
rect 10 942 50 944
rect 292 936 332 938
rect 10 924 50 926
rect 10 916 50 918
rect 292 918 332 920
rect 292 910 332 912
rect 292 892 332 894
rect 292 884 332 886
rect 10 880 50 882
rect 10 862 50 864
rect 10 854 50 856
rect 10 819 50 821
rect 10 811 50 813
rect 10 674 50 676
rect 10 666 50 668
rect 10 648 50 650
rect 10 640 50 642
rect 247 611 287 613
rect 10 604 50 606
rect 247 603 287 605
rect 10 586 50 588
rect 247 585 287 587
rect 10 578 50 580
rect 247 577 287 579
rect 10 543 50 545
rect 10 535 50 537
rect 10 388 50 390
rect 10 370 50 372
rect 10 362 50 364
rect 212 357 252 359
rect 212 339 252 341
rect 212 331 252 333
rect 10 320 50 322
rect 10 312 50 314
rect 11 177 51 179
rect 11 169 51 171
rect 185 158 225 160
rect 185 150 225 152
<< ndiffusion >>
rect 72 1058 172 1059
rect 72 1055 172 1056
rect 72 1040 172 1041
rect 72 1037 172 1038
rect 72 1032 172 1033
rect 72 1029 172 1030
rect 72 1014 172 1015
rect 72 1011 172 1012
rect 72 1006 172 1007
rect 72 1003 172 1004
rect 72 952 152 953
rect 72 949 152 950
rect 72 944 152 945
rect 72 941 152 942
rect 354 938 454 939
rect 354 935 454 936
rect 72 926 152 927
rect 72 923 152 924
rect 72 918 152 919
rect 354 920 454 921
rect 72 915 152 916
rect 354 917 454 918
rect 354 912 454 913
rect 354 909 454 910
rect 354 894 454 895
rect 354 891 454 892
rect 354 886 454 887
rect 72 882 132 883
rect 72 879 132 880
rect 354 883 454 884
rect 72 864 132 865
rect 72 861 132 862
rect 72 856 132 857
rect 72 853 132 854
rect 72 821 112 822
rect 72 818 112 819
rect 72 813 112 814
rect 72 810 112 811
rect 72 676 152 677
rect 72 673 152 674
rect 72 668 152 669
rect 72 665 152 666
rect 72 650 152 651
rect 72 647 152 648
rect 72 642 152 643
rect 72 639 152 640
rect 309 613 389 614
rect 72 606 132 607
rect 72 603 132 604
rect 309 610 389 611
rect 309 605 389 606
rect 309 602 389 603
rect 72 588 132 589
rect 72 585 132 586
rect 309 587 389 588
rect 72 580 132 581
rect 72 577 132 578
rect 309 584 389 585
rect 309 579 389 580
rect 309 576 389 577
rect 72 545 112 546
rect 72 542 112 543
rect 72 537 112 538
rect 72 534 112 535
rect 72 390 132 391
rect 72 387 132 388
rect 72 372 132 373
rect 72 369 132 370
rect 72 364 132 365
rect 72 361 132 362
rect 274 359 334 360
rect 274 356 334 357
rect 274 341 334 342
rect 274 338 334 339
rect 274 333 334 334
rect 274 330 334 331
rect 72 322 112 323
rect 72 319 112 320
rect 72 314 112 315
rect 72 311 112 312
rect 73 179 113 180
rect 73 176 113 177
rect 73 171 113 172
rect 73 168 113 169
rect 247 160 287 161
rect 247 157 287 158
rect 247 152 287 153
rect 247 149 287 150
<< pdiffusion >>
rect 10 1058 50 1059
rect 10 1055 50 1056
rect 10 1040 50 1041
rect 10 1037 50 1038
rect 10 1032 50 1033
rect 10 1029 50 1030
rect 10 1014 50 1015
rect 10 1011 50 1012
rect 10 1006 50 1007
rect 10 1003 50 1004
rect 10 952 50 953
rect 10 949 50 950
rect 10 944 50 945
rect 10 941 50 942
rect 292 938 332 939
rect 292 935 332 936
rect 10 926 50 927
rect 10 923 50 924
rect 10 918 50 919
rect 292 920 332 921
rect 292 917 332 918
rect 10 915 50 916
rect 292 912 332 913
rect 292 909 332 910
rect 292 894 332 895
rect 292 891 332 892
rect 10 882 50 883
rect 292 886 332 887
rect 292 883 332 884
rect 10 879 50 880
rect 10 864 50 865
rect 10 861 50 862
rect 10 856 50 857
rect 10 853 50 854
rect 10 821 50 822
rect 10 818 50 819
rect 10 813 50 814
rect 10 810 50 811
rect 10 676 50 677
rect 10 673 50 674
rect 10 668 50 669
rect 10 665 50 666
rect 10 650 50 651
rect 10 647 50 648
rect 10 642 50 643
rect 10 639 50 640
rect 10 606 50 607
rect 247 613 287 614
rect 247 610 287 611
rect 10 603 50 604
rect 247 605 287 606
rect 247 602 287 603
rect 10 588 50 589
rect 10 585 50 586
rect 10 580 50 581
rect 247 587 287 588
rect 247 584 287 585
rect 10 577 50 578
rect 247 579 287 580
rect 247 576 287 577
rect 10 545 50 546
rect 10 542 50 543
rect 10 537 50 538
rect 10 534 50 535
rect 10 390 50 391
rect 10 387 50 388
rect 10 372 50 373
rect 10 369 50 370
rect 10 364 50 365
rect 10 361 50 362
rect 212 359 252 360
rect 212 356 252 357
rect 212 341 252 342
rect 212 338 252 339
rect 212 333 252 334
rect 212 330 252 331
rect 10 322 50 323
rect 10 319 50 320
rect 10 314 50 315
rect 10 311 50 312
rect 11 179 51 180
rect 11 176 51 177
rect 11 171 51 172
rect 11 168 51 169
rect 185 160 225 161
rect 185 157 225 158
rect 185 152 225 153
rect 185 149 225 150
<< ndcontact >>
rect 72 1059 172 1063
rect 72 1051 172 1055
rect 72 1041 172 1045
rect 72 1033 172 1037
rect 72 1025 172 1029
rect 72 1015 172 1019
rect 72 1007 172 1011
rect 72 999 172 1003
rect 72 953 152 957
rect 72 945 152 949
rect 72 937 152 941
rect 354 939 454 943
rect 354 931 454 935
rect 72 927 152 931
rect 72 919 152 923
rect 354 921 454 925
rect 72 911 152 915
rect 354 913 454 917
rect 354 905 454 909
rect 354 895 454 899
rect 72 883 132 887
rect 354 887 454 891
rect 354 879 454 883
rect 72 875 132 879
rect 72 865 132 869
rect 72 857 132 861
rect 72 849 132 853
rect 72 822 112 826
rect 72 814 112 818
rect 72 806 112 810
rect 72 677 152 681
rect 72 669 152 673
rect 72 661 152 665
rect 72 651 152 655
rect 72 643 152 647
rect 72 635 152 639
rect 72 607 132 611
rect 309 614 389 618
rect 72 599 132 603
rect 309 606 389 610
rect 309 598 389 602
rect 72 589 132 593
rect 72 581 132 585
rect 309 588 389 592
rect 72 573 132 577
rect 309 580 389 584
rect 309 572 389 576
rect 72 546 112 550
rect 72 538 112 542
rect 72 530 112 534
rect 72 391 132 395
rect 72 383 132 387
rect 72 373 132 377
rect 72 365 132 369
rect 72 357 132 361
rect 274 360 334 364
rect 274 352 334 356
rect 274 342 334 346
rect 274 334 334 338
rect 72 323 112 327
rect 274 326 334 330
rect 72 315 112 319
rect 72 307 112 311
rect 73 180 113 184
rect 73 172 113 176
rect 73 164 113 168
rect 247 161 287 165
rect 247 153 287 157
rect 247 145 287 149
<< pdcontact >>
rect 10 1059 50 1063
rect 10 1051 50 1055
rect 10 1041 50 1045
rect 10 1033 50 1037
rect 10 1025 50 1029
rect 10 1015 50 1019
rect 10 1007 50 1011
rect 10 999 50 1003
rect 10 953 50 957
rect 10 945 50 949
rect 10 937 50 941
rect 292 939 332 943
rect 292 931 332 935
rect 10 927 50 931
rect 10 919 50 923
rect 292 921 332 925
rect 10 911 50 915
rect 292 913 332 917
rect 292 905 332 909
rect 292 895 332 899
rect 292 887 332 891
rect 10 883 50 887
rect 10 875 50 879
rect 292 879 332 883
rect 10 865 50 869
rect 10 857 50 861
rect 10 849 50 853
rect 10 822 50 826
rect 10 814 50 818
rect 10 806 50 810
rect 10 677 50 681
rect 10 669 50 673
rect 10 661 50 665
rect 10 651 50 655
rect 10 643 50 647
rect 10 635 50 639
rect 247 614 287 618
rect 10 607 50 611
rect 247 606 287 610
rect 10 599 50 603
rect 247 598 287 602
rect 10 589 50 593
rect 247 588 287 592
rect 10 581 50 585
rect 247 580 287 584
rect 10 573 50 577
rect 247 572 287 576
rect 10 546 50 550
rect 10 538 50 542
rect 10 530 50 534
rect 10 391 50 395
rect 10 383 50 387
rect 10 373 50 377
rect 10 365 50 369
rect 10 357 50 361
rect 212 360 252 364
rect 212 352 252 356
rect 212 342 252 346
rect 212 334 252 338
rect 10 323 50 327
rect 212 326 252 330
rect 10 315 50 319
rect 10 307 50 311
rect 11 180 51 184
rect 11 172 51 176
rect 11 164 51 168
rect 185 161 225 165
rect 185 153 225 157
rect 185 145 225 149
<< polysilicon >>
rect -3 1056 10 1058
rect 50 1056 72 1058
rect 172 1056 175 1058
rect -3 1038 10 1040
rect 50 1038 72 1040
rect 172 1038 175 1040
rect -3 1030 10 1032
rect 50 1030 72 1032
rect 172 1030 175 1032
rect -3 1012 10 1014
rect 50 1012 72 1014
rect 172 1012 175 1014
rect -3 1004 10 1006
rect 50 1004 72 1006
rect 172 1004 175 1006
rect -3 950 10 952
rect 50 950 72 952
rect 152 950 155 952
rect -3 942 10 944
rect 50 942 72 944
rect 152 942 155 944
rect 279 936 292 938
rect 332 936 354 938
rect 454 936 457 938
rect -3 924 10 926
rect 50 924 72 926
rect 152 924 155 926
rect -3 916 10 918
rect 50 916 72 918
rect 152 916 155 918
rect 279 918 292 920
rect 332 918 354 920
rect 454 918 457 920
rect 279 910 292 912
rect 332 910 354 912
rect 454 910 457 912
rect 279 892 292 894
rect 332 892 354 894
rect 454 892 457 894
rect 279 884 292 886
rect 332 884 354 886
rect 454 884 457 886
rect -3 880 10 882
rect 50 880 72 882
rect 132 880 135 882
rect -3 862 10 864
rect 50 862 72 864
rect 132 862 135 864
rect -3 854 10 856
rect 50 854 72 856
rect 132 854 135 856
rect -3 819 10 821
rect 50 819 72 821
rect 112 819 115 821
rect -3 811 10 813
rect 50 811 72 813
rect 112 811 115 813
rect -3 674 10 676
rect 50 674 72 676
rect 152 674 155 676
rect -3 666 10 668
rect 50 666 72 668
rect 152 666 155 668
rect -3 648 10 650
rect 50 648 72 650
rect 152 648 155 650
rect -3 640 10 642
rect 50 640 72 642
rect 152 640 155 642
rect 234 611 247 613
rect 287 611 309 613
rect 389 611 392 613
rect -3 604 10 606
rect 50 604 72 606
rect 132 604 135 606
rect 234 603 247 605
rect 287 603 309 605
rect 389 603 392 605
rect -3 586 10 588
rect 50 586 72 588
rect 132 586 135 588
rect 234 585 247 587
rect 287 585 309 587
rect 389 585 392 587
rect -3 578 10 580
rect 50 578 72 580
rect 132 578 135 580
rect 234 577 247 579
rect 287 577 309 579
rect 389 577 392 579
rect -3 543 10 545
rect 50 543 72 545
rect 112 543 115 545
rect -3 535 10 537
rect 50 535 72 537
rect 112 535 115 537
rect -3 388 10 390
rect 50 388 72 390
rect 132 388 135 390
rect -3 370 10 372
rect 50 370 72 372
rect 132 370 135 372
rect -3 362 10 364
rect 50 362 72 364
rect 132 362 135 364
rect 199 357 212 359
rect 252 357 274 359
rect 334 357 337 359
rect 199 339 212 341
rect 252 339 274 341
rect 334 339 337 341
rect 199 331 212 333
rect 252 331 274 333
rect 334 331 337 333
rect -3 320 10 322
rect 50 320 72 322
rect 112 320 115 322
rect -3 312 10 314
rect 50 312 72 314
rect 112 312 115 314
rect -2 177 11 179
rect 51 177 73 179
rect 113 177 116 179
rect -2 169 11 171
rect 51 169 73 171
rect 113 169 116 171
rect 172 158 185 160
rect 225 158 247 160
rect 287 158 290 160
rect 172 150 185 152
rect 225 150 247 152
rect 287 150 290 152
<< polycontact >>
rect -7 1055 -3 1059
rect -7 1037 -3 1041
rect -7 1029 -3 1033
rect -7 1011 -3 1015
rect -7 1003 -3 1007
rect -7 949 -3 953
rect -7 941 -3 945
rect 275 935 279 939
rect -7 923 -3 927
rect -7 915 -3 919
rect 275 917 279 921
rect 275 909 279 913
rect 275 891 279 895
rect -7 879 -3 883
rect 275 883 279 887
rect -7 861 -3 865
rect -7 853 -3 857
rect -7 818 -3 822
rect -7 810 -3 814
rect -7 673 -3 677
rect -7 665 -3 669
rect -7 647 -3 651
rect -7 639 -3 643
rect -7 603 -3 607
rect 230 610 234 614
rect 230 602 234 606
rect -7 585 -3 589
rect -7 577 -3 581
rect 230 584 234 588
rect 230 576 234 580
rect -7 542 -3 546
rect -7 534 -3 538
rect -7 387 -3 391
rect -7 369 -3 373
rect -7 361 -3 365
rect 195 356 199 360
rect 195 338 199 342
rect 195 330 199 334
rect -7 319 -3 323
rect -7 311 -3 315
rect -6 176 -2 180
rect -6 168 -2 172
rect 168 157 172 161
rect 168 149 172 153
<< metal1 >>
rect -12 1055 -7 1059
rect 2 1055 6 1080
rect 50 1059 58 1063
rect 172 1059 180 1063
rect 1 1051 10 1055
rect -12 1037 -7 1041
rect 2 1037 6 1051
rect 54 1045 58 1059
rect 50 1041 58 1045
rect 66 1051 72 1055
rect 66 1045 70 1051
rect 66 1041 72 1045
rect 1 1033 10 1037
rect -12 1029 -7 1033
rect -12 1011 -7 1015
rect 2 1011 6 1033
rect 54 1029 58 1041
rect 50 1025 59 1029
rect 66 1025 72 1029
rect 54 1019 58 1025
rect 50 1015 58 1019
rect 66 1019 70 1025
rect 66 1015 72 1019
rect 1 1007 10 1011
rect -12 1003 -7 1007
rect -11 949 -7 953
rect 2 949 6 1007
rect 54 1003 58 1015
rect 50 999 72 1003
rect 62 987 66 999
rect 62 983 269 987
rect 50 953 58 957
rect 152 953 160 957
rect 1 945 10 949
rect -11 941 -7 945
rect -12 923 -7 927
rect 2 923 6 945
rect 54 941 58 953
rect 50 937 59 941
rect 66 937 72 941
rect 265 939 269 983
rect 54 931 58 937
rect 50 927 58 931
rect 66 931 70 937
rect 265 935 275 939
rect 282 935 286 952
rect 332 939 340 943
rect 454 939 462 943
rect 265 934 269 935
rect 282 931 292 935
rect 66 927 72 931
rect 1 919 10 923
rect -12 915 -7 919
rect 2 887 6 919
rect 54 915 58 927
rect 177 917 275 921
rect 282 917 286 931
rect 336 925 340 939
rect 332 921 340 925
rect 348 931 354 935
rect 348 925 352 931
rect 348 921 354 925
rect 50 911 72 915
rect 62 906 66 911
rect 177 906 181 917
rect 282 913 292 917
rect 62 902 181 906
rect 196 909 275 913
rect 1 883 10 887
rect 132 883 139 887
rect -11 879 -7 883
rect -12 861 -7 865
rect 2 861 6 883
rect 50 875 58 879
rect 54 869 58 875
rect 50 865 58 869
rect 66 875 72 879
rect 66 869 70 875
rect 66 865 72 869
rect 1 857 10 861
rect -12 853 -7 857
rect -11 818 -7 822
rect 2 818 6 857
rect 54 853 58 865
rect 50 849 72 853
rect 65 844 69 849
rect 196 844 200 909
rect 65 840 200 844
rect 209 891 275 895
rect 282 891 286 913
rect 336 909 340 921
rect 332 905 341 909
rect 348 905 354 909
rect 336 899 340 905
rect 332 895 340 899
rect 348 899 352 905
rect 348 895 354 899
rect 50 822 58 826
rect 112 822 120 826
rect 1 814 10 818
rect -11 810 -7 814
rect 2 786 6 814
rect 54 810 58 822
rect 50 806 72 810
rect 65 801 69 806
rect 209 801 213 891
rect 282 887 292 891
rect 271 883 275 887
rect 65 797 213 801
rect 282 786 286 887
rect 336 883 340 895
rect 332 879 354 883
rect 344 837 348 879
rect 344 833 540 837
rect 536 826 540 833
rect 2 782 286 786
rect -35 673 -7 677
rect 2 673 6 782
rect 50 677 58 681
rect 152 677 160 681
rect 1 669 10 673
rect -29 665 -7 669
rect -21 647 -7 651
rect 2 647 6 669
rect 54 665 58 677
rect 50 661 59 665
rect 66 661 72 665
rect 54 655 58 661
rect 50 651 58 655
rect 66 655 70 661
rect 66 651 72 655
rect 1 643 10 647
rect -13 639 -7 643
rect 2 611 6 643
rect 54 639 58 651
rect 50 635 72 639
rect 62 622 66 635
rect 62 618 164 622
rect 160 614 164 618
rect 1 607 10 611
rect 132 607 139 611
rect 160 610 230 614
rect 238 610 242 624
rect 287 614 295 618
rect 389 614 397 618
rect -29 603 -7 607
rect -21 585 -7 589
rect 2 585 6 607
rect 238 606 247 610
rect 50 599 58 603
rect 54 593 58 599
rect 50 589 58 593
rect 66 599 72 603
rect 157 602 230 606
rect 66 593 70 599
rect 66 589 72 593
rect 1 581 10 585
rect -14 577 -7 581
rect -21 542 -7 546
rect 2 542 6 581
rect 54 577 58 589
rect 50 573 72 577
rect 64 569 68 573
rect 157 569 161 602
rect 64 565 161 569
rect 171 584 230 588
rect 238 584 242 606
rect 291 602 295 614
rect 287 598 296 602
rect 303 598 309 602
rect 291 592 295 598
rect 287 588 295 592
rect 303 592 307 598
rect 303 588 309 592
rect 50 546 58 550
rect 112 546 120 550
rect 1 538 10 542
rect -13 534 -7 538
rect 2 505 6 538
rect 54 534 58 546
rect 50 530 72 534
rect 61 526 65 530
rect 171 526 175 584
rect 238 580 247 584
rect 224 576 230 580
rect 61 522 175 526
rect 238 505 242 580
rect 291 576 295 588
rect 287 572 309 576
rect 296 524 300 572
rect 296 520 497 524
rect 2 501 242 505
rect 2 395 6 501
rect 1 391 10 395
rect 132 391 139 395
rect -29 387 -7 391
rect -21 369 -7 373
rect 2 369 6 391
rect 50 383 58 387
rect 54 377 58 383
rect 50 373 58 377
rect 66 383 72 387
rect 66 377 70 383
rect 66 373 72 377
rect 1 365 10 369
rect -13 361 -7 365
rect -24 319 -7 323
rect 2 319 6 365
rect 54 361 58 373
rect 202 364 206 376
rect 50 357 72 361
rect 202 360 212 364
rect 334 360 341 364
rect 62 349 66 357
rect 158 356 195 360
rect 158 349 162 356
rect 62 345 162 349
rect 170 338 195 342
rect 202 338 206 360
rect 252 352 260 356
rect 256 346 260 352
rect 252 342 260 346
rect 268 352 274 356
rect 268 346 272 352
rect 268 342 274 346
rect 50 323 58 327
rect 112 323 120 327
rect 1 315 10 319
rect -29 311 -7 315
rect 2 286 6 315
rect 54 311 58 323
rect 50 307 72 311
rect 63 302 67 307
rect 170 302 174 338
rect 202 334 212 338
rect 189 330 195 334
rect 63 298 174 302
rect 202 286 206 334
rect 256 330 260 342
rect 252 326 274 330
rect 264 304 268 326
rect 264 300 376 304
rect 2 282 206 286
rect -29 176 -6 180
rect 2 176 6 282
rect 51 180 59 184
rect 113 180 121 184
rect 2 172 11 176
rect -12 168 -6 172
rect 2 158 6 172
rect 55 168 59 180
rect 51 164 73 168
rect 64 161 68 164
rect 225 161 233 165
rect 287 161 295 165
rect 64 157 168 161
rect 176 153 185 157
rect 162 149 168 153
rect 229 149 233 161
rect 225 145 247 149
rect 236 132 240 145
rect 236 128 354 132
<< labels >>
rlabel metal1 162 149 165 153 1 g1
rlabel metal1 190 330 193 334 1 g2
rlabel metal1 225 576 228 580 1 g3
rlabel metal1 271 883 274 887 1 g4
rlabel metal1 -11 168 -8 172 1 g0
rlabel metal1 -12 1003 -9 1007 1 g0
rlabel metal1 -12 915 -9 919 1 g1
rlabel metal1 -12 853 -9 857 1 g2
rlabel metal1 -11 810 -8 814 1 g3
rlabel metal1 -12 639 -9 643 1 g0
rlabel metal1 -11 577 -8 581 1 g1
rlabel metal1 -11 534 -8 538 1 g2
rlabel metal1 -11 311 -8 315 1 g1
rlabel metal1 -11 176 -8 180 1 p1
rlabel metal1 -11 319 -8 323 1 p2
rlabel metal1 -11 542 -8 546 1 p3
rlabel metal1 -11 585 -8 589 1 p2
rlabel metal1 -11 603 -8 607 1 p3
rlabel metal1 -12 647 -9 651 1 p1
rlabel metal1 -12 665 -9 669 1 p2
rlabel metal1 -12 673 -9 677 1 p3
rlabel metal1 -11 818 -8 822 1 p4
rlabel metal1 -12 861 -9 865 1 p3
rlabel metal1 -11 879 -8 883 1 p4
rlabel metal1 -12 923 -9 927 1 p2
rlabel metal1 -11 941 -8 945 1 p3
rlabel metal1 -11 949 -8 953 1 p4
rlabel metal1 349 128 353 132 1 c2
rlabel metal1 370 300 374 304 1 c3
rlabel metal1 483 520 487 524 1 c4
rlabel metal1 527 833 531 837 1 c5
rlabel metal1 -12 1029 -9 1033 1 p2
rlabel metal1 -12 1011 -9 1015 1 p1
rlabel metal1 -12 1037 -9 1041 1 p3
rlabel metal1 -12 1055 -9 1059 1 p4
rlabel metal1 -11 361 -8 365 1 g0
rlabel metal1 -11 369 -8 373 1 p1
rlabel metal1 -12 387 -9 391 1 p2
<< end >>
